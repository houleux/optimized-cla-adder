magic
tech scmos
timestamp 1733175357
<< nwell >>
rect 1193 89 1587 127
rect 1745 125 1783 519
rect 1941 125 1979 519
rect 2969 284 3339 322
rect 2969 83 3348 121
rect 1193 -94 1587 -56
rect 1701 -100 1741 -38
rect 1789 -100 1829 -38
rect 1878 -100 1918 -38
rect 1966 -100 2006 -38
rect 1691 -147 1729 -106
rect 1779 -147 1817 -106
rect 1868 -147 1906 -106
rect 1956 -147 1994 -106
rect 2091 -151 2123 -86
rect 2202 -115 2234 -25
rect 2461 -35 2523 5
rect 2529 -23 2570 15
rect 2172 -151 2234 -115
rect 2340 -151 2372 -103
rect 2461 -221 2523 -181
rect 2529 -209 2570 -171
rect 2968 -198 3345 -160
rect 1188 -332 1582 -294
rect 1692 -362 1954 -330
rect 1967 -417 1999 -303
rect 2461 -436 2523 -396
rect 2529 -424 2570 -386
rect 2969 -462 3343 -424
rect 1188 -528 1582 -490
rect 1723 -893 1761 -499
rect 1919 -893 1957 -499
rect 2969 -663 3342 -625
<< ntransistor >>
rect 1789 427 1799 429
rect 1925 427 1935 429
rect 1789 356 1799 358
rect 1925 356 1935 358
rect 1789 320 1799 322
rect 1925 320 1935 322
rect 3059 268 3061 278
rect 1789 248 1799 250
rect 1925 248 1935 250
rect 3130 268 3132 278
rect 3166 268 3168 278
rect 3238 268 3240 278
rect 3274 268 3276 278
rect 3310 268 3312 278
rect 3326 268 3328 278
rect 1789 212 1799 214
rect 1925 212 1935 214
rect 1789 176 1799 178
rect 1925 176 1935 178
rect 1789 158 1799 160
rect 1925 158 1935 160
rect 1789 142 1799 144
rect 1925 142 1935 144
rect 1283 73 1285 83
rect 1354 73 1356 83
rect 1390 73 1392 83
rect 3059 127 3061 137
rect 3130 127 3132 137
rect 3166 127 3168 137
rect 1462 73 1464 83
rect 1498 73 1500 83
rect 1534 73 1536 83
rect 1552 73 1554 83
rect 1568 73 1570 83
rect 3238 127 3240 137
rect 3274 127 3276 137
rect 3310 127 3312 137
rect 3329 127 3331 137
rect 1283 -50 1285 -40
rect 1354 -50 1356 -40
rect 1390 -50 1392 -40
rect 1462 -50 1464 -40
rect 1498 -50 1500 -40
rect 1534 -50 1536 -40
rect 1552 -50 1554 -40
rect 1568 -50 1570 -40
rect 1747 -42 1757 -40
rect 1835 -42 1845 -40
rect 1924 -42 1934 -40
rect 2262 -38 2282 -36
rect 2012 -42 2022 -40
rect 2262 -50 2282 -48
rect 2463 -51 2465 -41
rect 2541 -42 2543 -32
rect 2557 -42 2559 -32
rect 2252 -68 2282 -66
rect 2252 -80 2282 -78
rect 2252 -92 2282 -90
rect 2042 -99 2062 -97
rect 2042 -111 2062 -109
rect 1738 -120 1748 -118
rect 1826 -120 1836 -118
rect 1915 -120 1925 -118
rect 2252 -116 2282 -114
rect 2293 -116 2323 -114
rect 2003 -120 2013 -118
rect 2042 -128 2062 -126
rect 2140 -128 2160 -126
rect 2252 -128 2282 -126
rect 2293 -128 2323 -126
rect 1738 -136 1748 -134
rect 1826 -136 1836 -134
rect 1915 -136 1925 -134
rect 2003 -136 2013 -134
rect 2042 -140 2062 -138
rect 2140 -140 2160 -138
rect 2252 -140 2282 -138
rect 2293 -140 2323 -138
rect 3058 -154 3060 -144
rect 3129 -154 3131 -144
rect 3165 -154 3167 -144
rect 3237 -154 3239 -144
rect 3273 -154 3275 -144
rect 3309 -154 3311 -144
rect 3326 -154 3328 -144
rect 2463 -237 2465 -227
rect 2541 -228 2543 -218
rect 2557 -228 2559 -218
rect 1278 -348 1280 -338
rect 1349 -348 1351 -338
rect 1385 -348 1387 -338
rect 1703 -310 1705 -290
rect 1715 -310 1717 -290
rect 1759 -310 1761 -290
rect 1771 -310 1773 -290
rect 1739 -321 1741 -311
rect 1812 -310 1814 -290
rect 1824 -310 1826 -290
rect 1795 -321 1797 -311
rect 1868 -310 1870 -290
rect 1880 -310 1882 -290
rect 1847 -321 1849 -311
rect 1903 -321 1905 -311
rect 1923 -321 1925 -311
rect 1941 -321 1943 -311
rect 2031 -316 2071 -314
rect 2031 -328 2071 -326
rect 1457 -348 1459 -338
rect 1493 -348 1495 -338
rect 1529 -348 1531 -338
rect 1547 -348 1549 -338
rect 1563 -348 1565 -338
rect 2031 -340 2071 -338
rect 2031 -352 2071 -350
rect 2031 -370 2071 -368
rect 2031 -382 2071 -380
rect 2031 -394 2071 -392
rect 2031 -406 2071 -404
rect 2463 -452 2465 -442
rect 2541 -443 2543 -433
rect 2557 -443 2559 -433
rect 1278 -484 1280 -474
rect 1349 -484 1351 -474
rect 1385 -484 1387 -474
rect 1457 -484 1459 -474
rect 1493 -484 1495 -474
rect 1529 -484 1531 -474
rect 1547 -484 1549 -474
rect 1563 -484 1565 -474
rect 3059 -478 3061 -468
rect 3130 -478 3132 -468
rect 3166 -478 3168 -468
rect 3238 -478 3240 -468
rect 3274 -478 3276 -468
rect 3310 -478 3312 -468
rect 3326 -478 3328 -468
rect 1767 -518 1777 -516
rect 1903 -518 1913 -516
rect 1767 -534 1777 -532
rect 1903 -534 1913 -532
rect 1767 -552 1777 -550
rect 1903 -552 1913 -550
rect 1767 -588 1777 -586
rect 1903 -588 1913 -586
rect 1767 -624 1777 -622
rect 1903 -624 1913 -622
rect 3059 -619 3061 -609
rect 3130 -619 3132 -609
rect 3166 -619 3168 -609
rect 3238 -619 3240 -609
rect 3274 -619 3276 -609
rect 3310 -619 3312 -609
rect 3326 -619 3328 -609
rect 1767 -696 1777 -694
rect 1903 -696 1913 -694
rect 1767 -732 1777 -730
rect 1903 -732 1913 -730
rect 1767 -803 1777 -801
rect 1903 -803 1913 -801
<< ptransistor >>
rect 1756 500 1776 502
rect 1948 500 1968 502
rect 1756 464 1776 466
rect 1948 464 1968 466
rect 1756 392 1776 394
rect 1948 392 1968 394
rect 2986 291 2988 311
rect 3022 291 3024 311
rect 1756 284 1776 286
rect 1948 284 1968 286
rect 3094 291 3096 311
rect 3202 291 3204 311
rect 3310 291 3312 311
rect 3326 291 3328 311
rect 1756 176 1776 178
rect 1948 176 1968 178
rect 1756 158 1776 160
rect 1948 158 1968 160
rect 1756 142 1776 144
rect 1948 142 1968 144
rect 1210 96 1212 116
rect 1246 96 1248 116
rect 1318 96 1320 116
rect 1426 96 1428 116
rect 1534 96 1536 116
rect 1552 96 1554 116
rect 1568 96 1570 116
rect 2986 94 2988 114
rect 3022 94 3024 114
rect 3094 94 3096 114
rect 3202 94 3204 114
rect 3310 94 3312 114
rect 3329 94 3331 114
rect 2467 -8 2517 -6
rect 2541 -17 2543 3
rect 2557 -17 2559 3
rect 1210 -83 1212 -63
rect 1246 -83 1248 -63
rect 1318 -83 1320 -63
rect 2467 -24 2517 -22
rect 1426 -83 1428 -63
rect 1534 -83 1536 -63
rect 1552 -83 1554 -63
rect 1568 -83 1570 -63
rect 1712 -94 1714 -44
rect 1728 -94 1730 -44
rect 1800 -94 1802 -44
rect 1816 -94 1818 -44
rect 1889 -94 1891 -44
rect 1905 -94 1907 -44
rect 2208 -38 2228 -36
rect 1977 -94 1979 -44
rect 1993 -94 1995 -44
rect 2208 -50 2228 -48
rect 2208 -68 2228 -66
rect 2208 -80 2228 -78
rect 2208 -92 2228 -90
rect 2097 -99 2117 -97
rect 2097 -111 2117 -109
rect 1703 -120 1723 -118
rect 1791 -120 1811 -118
rect 1880 -120 1900 -118
rect 1968 -120 1988 -118
rect 2208 -116 2228 -114
rect 2346 -116 2366 -114
rect 2097 -128 2117 -126
rect 2178 -128 2198 -126
rect 2208 -128 2228 -126
rect 2346 -128 2366 -126
rect 1703 -136 1723 -134
rect 1791 -136 1811 -134
rect 1880 -136 1900 -134
rect 1968 -136 1988 -134
rect 2097 -140 2117 -138
rect 2178 -140 2198 -138
rect 2208 -140 2228 -138
rect 2346 -140 2366 -138
rect 2467 -194 2517 -192
rect 2541 -203 2543 -183
rect 2557 -203 2559 -183
rect 2985 -187 2987 -167
rect 3021 -187 3023 -167
rect 3093 -187 3095 -167
rect 3201 -187 3203 -167
rect 2467 -210 2517 -208
rect 3309 -187 3311 -167
rect 3326 -187 3328 -167
rect 1205 -325 1207 -305
rect 1241 -325 1243 -305
rect 1313 -325 1315 -305
rect 1421 -325 1423 -305
rect 1529 -325 1531 -305
rect 1547 -325 1549 -305
rect 1563 -325 1565 -305
rect 1973 -316 1993 -314
rect 1973 -328 1993 -326
rect 1703 -356 1705 -336
rect 1715 -356 1717 -336
rect 1739 -356 1741 -336
rect 1759 -356 1761 -336
rect 1771 -356 1773 -336
rect 1795 -356 1797 -336
rect 1812 -356 1814 -336
rect 1824 -356 1826 -336
rect 1847 -356 1849 -336
rect 1868 -356 1870 -336
rect 1880 -356 1882 -336
rect 1903 -356 1905 -336
rect 1923 -356 1925 -336
rect 1941 -356 1943 -336
rect 1973 -340 1993 -338
rect 1973 -352 1993 -350
rect 1973 -370 1993 -368
rect 1973 -382 1993 -380
rect 1973 -394 1993 -392
rect 1973 -406 1993 -404
rect 2467 -409 2517 -407
rect 2541 -418 2543 -398
rect 2557 -418 2559 -398
rect 2467 -425 2517 -423
rect 1205 -517 1207 -497
rect 1241 -517 1243 -497
rect 1313 -517 1315 -497
rect 2986 -455 2988 -435
rect 3022 -455 3024 -435
rect 1421 -517 1423 -497
rect 3094 -455 3096 -435
rect 1529 -517 1531 -497
rect 1547 -517 1549 -497
rect 1563 -517 1565 -497
rect 3202 -455 3204 -435
rect 3310 -455 3312 -435
rect 3326 -455 3328 -435
rect 1734 -518 1754 -516
rect 1926 -518 1946 -516
rect 1734 -534 1754 -532
rect 1926 -534 1946 -532
rect 1734 -552 1754 -550
rect 1926 -552 1946 -550
rect 2986 -652 2988 -632
rect 3022 -652 3024 -632
rect 3094 -652 3096 -632
rect 1734 -660 1754 -658
rect 1926 -660 1946 -658
rect 3202 -652 3204 -632
rect 3310 -652 3312 -632
rect 3326 -652 3328 -632
rect 1734 -768 1754 -766
rect 1926 -768 1946 -766
rect 1734 -840 1754 -838
rect 1926 -840 1946 -838
rect 1734 -876 1754 -874
rect 1926 -876 1946 -874
<< ndiffusion >>
rect 1798 430 1799 434
rect 1789 429 1799 430
rect 1789 426 1799 427
rect 1925 430 1926 434
rect 1925 429 1935 430
rect 1925 426 1935 427
rect 1798 359 1799 363
rect 1789 358 1799 359
rect 1925 359 1926 363
rect 1925 358 1935 359
rect 1789 355 1799 356
rect 1798 351 1799 355
rect 1925 355 1935 356
rect 1925 351 1926 355
rect 1798 323 1799 327
rect 1789 322 1799 323
rect 1789 319 1799 320
rect 1925 323 1926 327
rect 1925 322 1935 323
rect 1925 319 1935 320
rect 1798 251 1799 255
rect 3058 269 3059 278
rect 3054 268 3059 269
rect 3061 268 3062 278
rect 1789 250 1799 251
rect 1789 247 1799 248
rect 1798 243 1799 247
rect 1925 251 1926 255
rect 1925 250 1935 251
rect 3129 269 3130 278
rect 3125 268 3130 269
rect 3132 269 3133 278
rect 3132 268 3137 269
rect 3165 269 3166 278
rect 3161 268 3166 269
rect 3168 268 3169 278
rect 1925 247 1935 248
rect 1925 243 1926 247
rect 3237 269 3238 278
rect 3233 268 3238 269
rect 3240 269 3241 278
rect 3240 268 3245 269
rect 3273 269 3274 278
rect 3269 268 3274 269
rect 3276 268 3277 278
rect 3309 268 3310 278
rect 3312 269 3313 278
rect 3312 268 3317 269
rect 3325 268 3326 278
rect 3328 269 3329 278
rect 3328 268 3333 269
rect 1798 215 1799 219
rect 1789 214 1799 215
rect 1925 215 1926 219
rect 1925 214 1935 215
rect 1789 211 1799 212
rect 1925 211 1935 212
rect 1789 178 1799 179
rect 1925 178 1935 179
rect 1789 175 1799 176
rect 1798 171 1799 175
rect 1925 175 1935 176
rect 1925 171 1926 175
rect 1789 160 1799 161
rect 1925 160 1935 161
rect 1789 157 1799 158
rect 1798 153 1799 157
rect 1925 157 1935 158
rect 1925 153 1926 157
rect 1789 144 1799 145
rect 1925 144 1935 145
rect 1282 74 1283 83
rect 1278 73 1283 74
rect 1285 73 1286 83
rect 1789 141 1799 142
rect 1798 137 1799 141
rect 1925 141 1935 142
rect 1925 137 1926 141
rect 1353 74 1354 83
rect 1349 73 1354 74
rect 1356 74 1357 83
rect 1356 73 1361 74
rect 1389 74 1390 83
rect 1385 73 1390 74
rect 1392 73 1393 83
rect 3054 136 3059 137
rect 3058 127 3059 136
rect 3061 127 3062 137
rect 3125 136 3130 137
rect 3129 127 3130 136
rect 3132 136 3137 137
rect 3132 127 3133 136
rect 3161 136 3166 137
rect 3165 127 3166 136
rect 3168 127 3169 137
rect 1461 74 1462 83
rect 1457 73 1462 74
rect 1464 74 1465 83
rect 1464 73 1469 74
rect 1497 74 1498 83
rect 1493 73 1498 74
rect 1500 73 1501 83
rect 1533 73 1534 83
rect 1536 74 1537 83
rect 1536 73 1541 74
rect 1551 73 1552 83
rect 1554 74 1555 83
rect 1554 73 1559 74
rect 1567 73 1568 83
rect 1570 74 1571 83
rect 3233 136 3238 137
rect 3237 127 3238 136
rect 3240 136 3245 137
rect 3240 127 3241 136
rect 3269 136 3274 137
rect 3273 127 3274 136
rect 3276 127 3277 137
rect 3309 127 3310 137
rect 3312 136 3317 137
rect 3312 127 3313 136
rect 3328 127 3329 137
rect 3331 136 3336 137
rect 3331 127 3332 136
rect 1570 73 1575 74
rect 1278 -41 1283 -40
rect 1282 -50 1283 -41
rect 1285 -50 1286 -40
rect 1349 -41 1354 -40
rect 1353 -50 1354 -41
rect 1356 -41 1361 -40
rect 1356 -50 1357 -41
rect 1385 -41 1390 -40
rect 1389 -50 1390 -41
rect 1392 -50 1393 -40
rect 1457 -41 1462 -40
rect 1461 -50 1462 -41
rect 1464 -41 1469 -40
rect 1464 -50 1465 -41
rect 1493 -41 1498 -40
rect 1497 -50 1498 -41
rect 1500 -50 1501 -40
rect 1533 -50 1534 -40
rect 1536 -41 1541 -40
rect 1536 -50 1537 -41
rect 1551 -50 1552 -40
rect 1554 -41 1559 -40
rect 1554 -50 1555 -41
rect 1567 -50 1568 -40
rect 1570 -41 1575 -40
rect 1570 -50 1571 -41
rect 1747 -40 1757 -39
rect 1747 -43 1757 -42
rect 1835 -40 1845 -39
rect 1835 -43 1845 -42
rect 1924 -40 1934 -39
rect 1924 -43 1934 -42
rect 2267 -35 2282 -31
rect 2262 -36 2282 -35
rect 2012 -40 2022 -39
rect 2012 -43 2022 -42
rect 2262 -48 2282 -38
rect 2262 -51 2282 -50
rect 2462 -51 2463 -41
rect 2465 -51 2466 -41
rect 2540 -42 2541 -32
rect 2543 -34 2548 -32
rect 2543 -42 2544 -34
rect 2556 -42 2557 -32
rect 2559 -34 2564 -32
rect 2559 -42 2560 -34
rect 2262 -55 2277 -51
rect 2257 -65 2282 -61
rect 2252 -66 2282 -65
rect 2252 -78 2282 -68
rect 2252 -90 2282 -80
rect 2042 -96 2057 -92
rect 2042 -97 2062 -96
rect 2252 -93 2282 -92
rect 2252 -97 2277 -93
rect 2042 -109 2062 -99
rect 2042 -112 2062 -111
rect 1738 -118 1748 -117
rect 1826 -118 1836 -117
rect 1915 -118 1925 -117
rect 2047 -116 2062 -112
rect 2257 -113 2282 -109
rect 2252 -114 2282 -113
rect 2293 -113 2318 -109
rect 2293 -114 2323 -113
rect 2003 -118 2013 -117
rect 1738 -121 1748 -120
rect 1738 -125 1740 -121
rect 1826 -121 1836 -120
rect 1826 -125 1828 -121
rect 1915 -121 1925 -120
rect 1915 -125 1917 -121
rect 2003 -121 2013 -120
rect 2003 -125 2005 -121
rect 2042 -125 2057 -121
rect 2042 -126 2062 -125
rect 2140 -125 2155 -121
rect 2140 -126 2160 -125
rect 2252 -126 2282 -116
rect 2293 -126 2323 -116
rect 1738 -134 1748 -133
rect 1826 -134 1836 -133
rect 1915 -134 1925 -133
rect 2003 -134 2013 -133
rect 1738 -137 1748 -136
rect 1738 -141 1740 -137
rect 1826 -137 1836 -136
rect 1826 -141 1828 -137
rect 1915 -137 1925 -136
rect 1915 -141 1917 -137
rect 2003 -137 2013 -136
rect 2003 -141 2005 -137
rect 2042 -138 2062 -128
rect 2140 -138 2160 -128
rect 2252 -138 2282 -128
rect 2293 -138 2323 -128
rect 2042 -141 2062 -140
rect 2047 -145 2062 -141
rect 2140 -141 2160 -140
rect 2145 -145 2160 -141
rect 2252 -141 2282 -140
rect 2252 -145 2277 -141
rect 2293 -141 2323 -140
rect 2298 -145 2323 -141
rect 3053 -145 3058 -144
rect 3057 -154 3058 -145
rect 3060 -154 3061 -144
rect 3124 -145 3129 -144
rect 3128 -154 3129 -145
rect 3131 -145 3136 -144
rect 3131 -154 3132 -145
rect 3160 -145 3165 -144
rect 3164 -154 3165 -145
rect 3167 -154 3168 -144
rect 3232 -145 3237 -144
rect 3236 -154 3237 -145
rect 3239 -145 3244 -144
rect 3239 -154 3240 -145
rect 3268 -145 3273 -144
rect 3272 -154 3273 -145
rect 3275 -154 3276 -144
rect 3308 -154 3309 -144
rect 3311 -145 3316 -144
rect 3311 -154 3312 -145
rect 3325 -154 3326 -144
rect 3328 -145 3333 -144
rect 3328 -154 3329 -145
rect 2462 -237 2463 -227
rect 2465 -237 2466 -227
rect 2540 -228 2541 -218
rect 2543 -220 2548 -218
rect 2543 -228 2544 -220
rect 2556 -228 2557 -218
rect 2559 -220 2564 -218
rect 2559 -228 2560 -220
rect 1277 -347 1278 -338
rect 1273 -348 1278 -347
rect 1280 -348 1281 -338
rect 1348 -347 1349 -338
rect 1344 -348 1349 -347
rect 1351 -347 1352 -338
rect 1351 -348 1356 -347
rect 1384 -347 1385 -338
rect 1380 -348 1385 -347
rect 1387 -348 1388 -338
rect 1702 -295 1703 -290
rect 1698 -310 1703 -295
rect 1705 -310 1715 -290
rect 1717 -305 1722 -290
rect 1758 -295 1759 -290
rect 1717 -310 1718 -305
rect 1754 -310 1759 -295
rect 1761 -310 1771 -290
rect 1773 -305 1778 -290
rect 1811 -295 1812 -290
rect 1773 -310 1774 -305
rect 1738 -315 1739 -311
rect 1734 -321 1739 -315
rect 1741 -315 1746 -311
rect 1741 -321 1742 -315
rect 1807 -310 1812 -295
rect 1814 -310 1824 -290
rect 1826 -305 1831 -290
rect 1867 -295 1868 -290
rect 1826 -310 1827 -305
rect 1794 -316 1795 -311
rect 1790 -321 1795 -316
rect 1797 -315 1802 -311
rect 1797 -321 1798 -315
rect 1863 -310 1868 -295
rect 1870 -310 1880 -290
rect 1882 -305 1887 -290
rect 1882 -310 1883 -305
rect 1846 -316 1847 -311
rect 1842 -321 1847 -316
rect 1849 -315 1854 -311
rect 1849 -321 1850 -315
rect 1902 -316 1903 -311
rect 1898 -321 1903 -316
rect 1905 -315 1910 -311
rect 1905 -321 1906 -315
rect 1922 -316 1923 -311
rect 1918 -321 1923 -316
rect 1925 -315 1930 -311
rect 1925 -321 1926 -315
rect 1940 -316 1941 -311
rect 1936 -321 1941 -316
rect 1943 -315 1948 -311
rect 2031 -313 2066 -309
rect 2031 -314 2071 -313
rect 1943 -321 1944 -315
rect 2031 -326 2071 -316
rect 1456 -347 1457 -338
rect 1452 -348 1457 -347
rect 1459 -347 1460 -338
rect 1459 -348 1464 -347
rect 1492 -347 1493 -338
rect 1488 -348 1493 -347
rect 1495 -348 1496 -338
rect 1528 -348 1529 -338
rect 1531 -347 1532 -338
rect 1531 -348 1536 -347
rect 1546 -348 1547 -338
rect 1549 -347 1550 -338
rect 1549 -348 1554 -347
rect 1562 -348 1563 -338
rect 1565 -347 1566 -338
rect 1565 -348 1570 -347
rect 2031 -338 2071 -328
rect 2031 -350 2071 -340
rect 2031 -353 2071 -352
rect 2036 -357 2071 -353
rect 2031 -367 2066 -363
rect 2031 -368 2071 -367
rect 2031 -380 2071 -370
rect 2031 -392 2071 -382
rect 2031 -404 2071 -394
rect 2031 -407 2071 -406
rect 2036 -411 2071 -407
rect 2462 -452 2463 -442
rect 2465 -452 2466 -442
rect 2540 -443 2541 -433
rect 2543 -435 2548 -433
rect 2543 -443 2544 -435
rect 2556 -443 2557 -433
rect 2559 -435 2564 -433
rect 2559 -443 2560 -435
rect 1273 -475 1278 -474
rect 1277 -484 1278 -475
rect 1280 -484 1281 -474
rect 1344 -475 1349 -474
rect 1348 -484 1349 -475
rect 1351 -475 1356 -474
rect 1351 -484 1352 -475
rect 1380 -475 1385 -474
rect 1384 -484 1385 -475
rect 1387 -484 1388 -474
rect 1452 -475 1457 -474
rect 1456 -484 1457 -475
rect 1459 -475 1464 -474
rect 1459 -484 1460 -475
rect 1488 -475 1493 -474
rect 1492 -484 1493 -475
rect 1495 -484 1496 -474
rect 1528 -484 1529 -474
rect 1531 -475 1536 -474
rect 1531 -484 1532 -475
rect 1546 -484 1547 -474
rect 1549 -475 1554 -474
rect 1549 -484 1550 -475
rect 1562 -484 1563 -474
rect 1565 -475 1570 -474
rect 1565 -484 1566 -475
rect 3058 -477 3059 -468
rect 3054 -478 3059 -477
rect 3061 -478 3062 -468
rect 3129 -477 3130 -468
rect 3125 -478 3130 -477
rect 3132 -477 3133 -468
rect 3132 -478 3137 -477
rect 3165 -477 3166 -468
rect 3161 -478 3166 -477
rect 3168 -478 3169 -468
rect 3237 -477 3238 -468
rect 3233 -478 3238 -477
rect 3240 -477 3241 -468
rect 3240 -478 3245 -477
rect 3273 -477 3274 -468
rect 3269 -478 3274 -477
rect 3276 -478 3277 -468
rect 3309 -478 3310 -468
rect 3312 -477 3313 -468
rect 3312 -478 3317 -477
rect 3325 -478 3326 -468
rect 3328 -477 3329 -468
rect 3328 -478 3333 -477
rect 1776 -515 1777 -511
rect 1767 -516 1777 -515
rect 1903 -515 1904 -511
rect 1903 -516 1913 -515
rect 1767 -519 1777 -518
rect 1903 -519 1913 -518
rect 1776 -531 1777 -527
rect 1767 -532 1777 -531
rect 1903 -531 1904 -527
rect 1903 -532 1913 -531
rect 1767 -535 1777 -534
rect 1903 -535 1913 -534
rect 1776 -549 1777 -545
rect 1767 -550 1777 -549
rect 1903 -549 1904 -545
rect 1903 -550 1913 -549
rect 1767 -553 1777 -552
rect 1903 -553 1913 -552
rect 1767 -586 1777 -585
rect 1903 -586 1913 -585
rect 1767 -589 1777 -588
rect 1776 -593 1777 -589
rect 1903 -589 1913 -588
rect 1903 -593 1904 -589
rect 1776 -621 1777 -617
rect 1767 -622 1777 -621
rect 1767 -625 1777 -624
rect 1776 -629 1777 -625
rect 1903 -621 1904 -617
rect 1903 -622 1913 -621
rect 1903 -625 1913 -624
rect 1903 -629 1904 -625
rect 3054 -610 3059 -609
rect 3058 -619 3059 -610
rect 3061 -619 3062 -609
rect 3125 -610 3130 -609
rect 3129 -619 3130 -610
rect 3132 -610 3137 -609
rect 3132 -619 3133 -610
rect 3161 -610 3166 -609
rect 3165 -619 3166 -610
rect 3168 -619 3169 -609
rect 3233 -610 3238 -609
rect 3237 -619 3238 -610
rect 3240 -610 3245 -609
rect 3240 -619 3241 -610
rect 3269 -610 3274 -609
rect 3273 -619 3274 -610
rect 3276 -619 3277 -609
rect 3309 -619 3310 -609
rect 3312 -610 3317 -609
rect 3312 -619 3313 -610
rect 3325 -619 3326 -609
rect 3328 -610 3333 -609
rect 3328 -619 3329 -610
rect 1767 -694 1777 -693
rect 1767 -697 1777 -696
rect 1776 -701 1777 -697
rect 1903 -694 1913 -693
rect 1903 -697 1913 -696
rect 1903 -701 1904 -697
rect 1776 -729 1777 -725
rect 1767 -730 1777 -729
rect 1903 -729 1904 -725
rect 1903 -730 1913 -729
rect 1767 -733 1777 -732
rect 1776 -737 1777 -733
rect 1903 -733 1913 -732
rect 1903 -737 1904 -733
rect 1767 -801 1777 -800
rect 1767 -804 1777 -803
rect 1776 -808 1777 -804
rect 1903 -801 1913 -800
rect 1903 -804 1913 -803
rect 1903 -808 1904 -804
<< pdiffusion >>
rect 1756 502 1776 503
rect 1948 502 1968 503
rect 1756 499 1776 500
rect 1948 499 1968 500
rect 1756 466 1776 467
rect 1948 466 1968 467
rect 1756 463 1776 464
rect 1948 463 1968 464
rect 1756 394 1776 395
rect 1756 391 1776 392
rect 1948 394 1968 395
rect 1948 391 1968 392
rect 1756 286 1776 287
rect 2985 291 2986 311
rect 2988 291 2989 311
rect 3021 291 3022 311
rect 3024 291 3025 311
rect 1948 286 1968 287
rect 1756 283 1776 284
rect 1948 283 1968 284
rect 3093 291 3094 311
rect 3096 291 3097 311
rect 3201 291 3202 311
rect 3204 291 3205 311
rect 3309 291 3310 311
rect 3312 291 3313 311
rect 3325 291 3326 311
rect 3328 291 3329 311
rect 1756 178 1776 179
rect 1948 178 1968 179
rect 1756 175 1776 176
rect 1948 175 1968 176
rect 1756 160 1776 161
rect 1948 160 1968 161
rect 1756 157 1776 158
rect 1948 157 1968 158
rect 1756 144 1776 145
rect 1948 144 1968 145
rect 1756 141 1776 142
rect 1209 96 1210 116
rect 1212 96 1213 116
rect 1245 96 1246 116
rect 1248 96 1249 116
rect 1317 96 1318 116
rect 1320 96 1321 116
rect 1948 141 1968 142
rect 1425 96 1426 116
rect 1428 96 1429 116
rect 1533 96 1534 116
rect 1536 96 1537 116
rect 1551 96 1552 116
rect 1554 96 1555 116
rect 1567 96 1568 116
rect 1570 96 1571 116
rect 2985 94 2986 114
rect 2988 94 2989 114
rect 3021 94 3022 114
rect 3024 94 3025 114
rect 3093 94 3094 114
rect 3096 94 3097 114
rect 3201 94 3202 114
rect 3204 94 3205 114
rect 3309 94 3310 114
rect 3312 94 3313 114
rect 3328 94 3329 114
rect 3331 94 3332 114
rect 2467 -6 2517 -5
rect 2467 -9 2517 -8
rect 2540 -17 2541 3
rect 2543 -17 2544 3
rect 2556 -17 2557 3
rect 2559 -17 2560 3
rect 1209 -83 1210 -63
rect 1212 -83 1213 -63
rect 1245 -83 1246 -63
rect 1248 -83 1249 -63
rect 1317 -83 1318 -63
rect 1320 -83 1321 -63
rect 2467 -22 2517 -21
rect 2467 -25 2517 -24
rect 1425 -83 1426 -63
rect 1428 -83 1429 -63
rect 1533 -83 1534 -63
rect 1536 -83 1537 -63
rect 1551 -83 1552 -63
rect 1554 -83 1555 -63
rect 1567 -83 1568 -63
rect 1570 -83 1571 -63
rect 1711 -94 1712 -44
rect 1714 -94 1715 -44
rect 1727 -94 1728 -44
rect 1730 -94 1731 -44
rect 1799 -94 1800 -44
rect 1802 -94 1803 -44
rect 1815 -94 1816 -44
rect 1818 -94 1819 -44
rect 2214 -35 2228 -31
rect 1888 -94 1889 -44
rect 1891 -94 1892 -44
rect 1904 -94 1905 -44
rect 1907 -94 1908 -44
rect 2208 -36 2228 -35
rect 2208 -41 2228 -38
rect 1976 -94 1977 -44
rect 1979 -94 1980 -44
rect 1992 -94 1993 -44
rect 1995 -94 1996 -44
rect 2208 -45 2222 -41
rect 2208 -48 2228 -45
rect 2208 -51 2228 -50
rect 2214 -55 2228 -51
rect 2208 -65 2222 -61
rect 2208 -66 2228 -65
rect 2208 -71 2228 -68
rect 2214 -75 2228 -71
rect 2208 -78 2228 -75
rect 2208 -83 2228 -80
rect 2208 -87 2222 -83
rect 2208 -90 2228 -87
rect 2097 -96 2111 -92
rect 2097 -97 2117 -96
rect 2208 -93 2228 -92
rect 2214 -97 2228 -93
rect 2097 -102 2117 -99
rect 2103 -106 2117 -102
rect 2097 -109 2117 -106
rect 1703 -118 1723 -117
rect 1791 -118 1811 -117
rect 1880 -118 1900 -117
rect 1968 -118 1988 -117
rect 2097 -112 2117 -111
rect 2097 -116 2111 -112
rect 2208 -113 2222 -109
rect 2208 -114 2228 -113
rect 2352 -113 2366 -109
rect 2346 -114 2366 -113
rect 2208 -119 2228 -116
rect 1703 -121 1723 -120
rect 1791 -121 1811 -120
rect 1880 -121 1900 -120
rect 1968 -121 1988 -120
rect 2097 -125 2111 -121
rect 2097 -126 2117 -125
rect 2178 -125 2192 -121
rect 2178 -126 2198 -125
rect 2214 -123 2228 -119
rect 2208 -126 2228 -123
rect 2346 -119 2366 -116
rect 2346 -123 2360 -119
rect 2346 -126 2366 -123
rect 1703 -134 1723 -133
rect 1791 -134 1811 -133
rect 1880 -134 1900 -133
rect 1968 -134 1988 -133
rect 1703 -137 1723 -136
rect 1791 -137 1811 -136
rect 1880 -137 1900 -136
rect 1968 -137 1988 -136
rect 2097 -131 2117 -128
rect 2103 -135 2117 -131
rect 2097 -138 2117 -135
rect 2178 -131 2198 -128
rect 2184 -135 2198 -131
rect 2178 -138 2198 -135
rect 2208 -131 2228 -128
rect 2208 -135 2222 -131
rect 2208 -138 2228 -135
rect 2346 -131 2366 -128
rect 2352 -135 2366 -131
rect 2346 -138 2366 -135
rect 2097 -141 2117 -140
rect 2097 -145 2111 -141
rect 2178 -141 2198 -140
rect 2178 -145 2192 -141
rect 2208 -141 2228 -140
rect 2214 -145 2228 -141
rect 2346 -141 2366 -140
rect 2346 -145 2360 -141
rect 2467 -192 2517 -191
rect 2467 -195 2517 -194
rect 2540 -203 2541 -183
rect 2543 -203 2544 -183
rect 2556 -203 2557 -183
rect 2559 -203 2560 -183
rect 2984 -187 2985 -167
rect 2987 -187 2988 -167
rect 3020 -187 3021 -167
rect 3023 -187 3024 -167
rect 3092 -187 3093 -167
rect 3095 -187 3096 -167
rect 3200 -187 3201 -167
rect 3203 -187 3204 -167
rect 2467 -208 2517 -207
rect 2467 -211 2517 -210
rect 3308 -187 3309 -167
rect 3311 -187 3312 -167
rect 3325 -187 3326 -167
rect 3328 -187 3329 -167
rect 1204 -325 1205 -305
rect 1207 -325 1208 -305
rect 1240 -325 1241 -305
rect 1243 -325 1244 -305
rect 1312 -325 1313 -305
rect 1315 -325 1316 -305
rect 1420 -325 1421 -305
rect 1423 -325 1424 -305
rect 1528 -325 1529 -305
rect 1531 -325 1532 -305
rect 1546 -325 1547 -305
rect 1549 -325 1550 -305
rect 1562 -325 1563 -305
rect 1565 -325 1566 -305
rect 1979 -313 1993 -309
rect 1973 -314 1993 -313
rect 1973 -319 1993 -316
rect 1973 -323 1987 -319
rect 1973 -326 1993 -323
rect 1973 -331 1993 -328
rect 1979 -335 1993 -331
rect 1698 -350 1703 -336
rect 1702 -356 1703 -350
rect 1705 -342 1708 -336
rect 1712 -342 1715 -336
rect 1705 -356 1715 -342
rect 1717 -350 1722 -336
rect 1717 -356 1718 -350
rect 1734 -350 1739 -336
rect 1738 -356 1739 -350
rect 1741 -342 1742 -336
rect 1741 -356 1746 -342
rect 1754 -350 1759 -336
rect 1758 -356 1759 -350
rect 1761 -342 1764 -336
rect 1768 -342 1771 -336
rect 1761 -356 1771 -342
rect 1773 -350 1778 -336
rect 1773 -356 1774 -350
rect 1790 -350 1795 -336
rect 1794 -356 1795 -350
rect 1797 -342 1798 -336
rect 1797 -356 1802 -342
rect 1807 -350 1812 -336
rect 1811 -356 1812 -350
rect 1814 -342 1817 -336
rect 1821 -342 1824 -336
rect 1814 -356 1824 -342
rect 1826 -350 1831 -336
rect 1826 -356 1827 -350
rect 1842 -350 1847 -336
rect 1846 -356 1847 -350
rect 1849 -342 1850 -336
rect 1849 -356 1854 -342
rect 1863 -350 1868 -336
rect 1867 -356 1868 -350
rect 1870 -342 1873 -336
rect 1877 -342 1880 -336
rect 1870 -356 1880 -342
rect 1882 -350 1887 -336
rect 1882 -356 1883 -350
rect 1898 -350 1903 -336
rect 1902 -356 1903 -350
rect 1905 -342 1906 -336
rect 1905 -356 1910 -342
rect 1918 -350 1923 -336
rect 1922 -356 1923 -350
rect 1925 -342 1926 -336
rect 1925 -356 1930 -342
rect 1936 -350 1941 -336
rect 1940 -356 1941 -350
rect 1943 -342 1944 -336
rect 1973 -338 1993 -335
rect 1943 -356 1948 -342
rect 1973 -343 1993 -340
rect 1973 -347 1987 -343
rect 1973 -350 1993 -347
rect 1973 -353 1993 -352
rect 1979 -357 1993 -353
rect 1979 -367 1993 -363
rect 1973 -368 1993 -367
rect 1973 -373 1993 -370
rect 1973 -377 1987 -373
rect 1973 -380 1993 -377
rect 1973 -385 1993 -382
rect 1979 -389 1993 -385
rect 1973 -392 1993 -389
rect 1973 -397 1993 -394
rect 1973 -401 1987 -397
rect 1973 -404 1993 -401
rect 1973 -407 1993 -406
rect 1979 -411 1993 -407
rect 2467 -407 2517 -406
rect 2467 -410 2517 -409
rect 2540 -418 2541 -398
rect 2543 -418 2544 -398
rect 2556 -418 2557 -398
rect 2559 -418 2560 -398
rect 2467 -423 2517 -422
rect 2467 -426 2517 -425
rect 1204 -517 1205 -497
rect 1207 -517 1208 -497
rect 1240 -517 1241 -497
rect 1243 -517 1244 -497
rect 1312 -517 1313 -497
rect 1315 -517 1316 -497
rect 2985 -455 2986 -435
rect 2988 -455 2989 -435
rect 3021 -455 3022 -435
rect 3024 -455 3025 -435
rect 1420 -517 1421 -497
rect 1423 -517 1424 -497
rect 3093 -455 3094 -435
rect 3096 -455 3097 -435
rect 1528 -517 1529 -497
rect 1531 -517 1532 -497
rect 1546 -517 1547 -497
rect 1549 -517 1550 -497
rect 1562 -517 1563 -497
rect 1565 -517 1566 -497
rect 3201 -455 3202 -435
rect 3204 -455 3205 -435
rect 3309 -455 3310 -435
rect 3312 -455 3313 -435
rect 3325 -455 3326 -435
rect 3328 -455 3329 -435
rect 1734 -516 1754 -515
rect 1926 -516 1946 -515
rect 1734 -519 1754 -518
rect 1926 -519 1946 -518
rect 1734 -532 1754 -531
rect 1926 -532 1946 -531
rect 1734 -535 1754 -534
rect 1926 -535 1946 -534
rect 1734 -550 1754 -549
rect 1926 -550 1946 -549
rect 1734 -553 1754 -552
rect 1926 -553 1946 -552
rect 2985 -652 2986 -632
rect 2988 -652 2989 -632
rect 3021 -652 3022 -632
rect 3024 -652 3025 -632
rect 1734 -658 1754 -657
rect 3093 -652 3094 -632
rect 3096 -652 3097 -632
rect 1926 -658 1946 -657
rect 1734 -661 1754 -660
rect 1926 -661 1946 -660
rect 3201 -652 3202 -632
rect 3204 -652 3205 -632
rect 3309 -652 3310 -632
rect 3312 -652 3313 -632
rect 3325 -652 3326 -632
rect 3328 -652 3329 -632
rect 1734 -766 1754 -765
rect 1734 -769 1754 -768
rect 1926 -766 1946 -765
rect 1926 -769 1946 -768
rect 1734 -838 1754 -837
rect 1926 -838 1946 -837
rect 1734 -841 1754 -840
rect 1926 -841 1946 -840
rect 1734 -874 1754 -873
rect 1926 -874 1946 -873
rect 1734 -877 1754 -876
rect 1926 -877 1946 -876
<< ndcontact >>
rect 1789 430 1798 434
rect 1789 422 1799 426
rect 1926 430 1935 434
rect 1925 422 1935 426
rect 1789 359 1798 363
rect 1926 359 1935 363
rect 1789 351 1798 355
rect 1926 351 1935 355
rect 1789 323 1798 327
rect 1789 315 1799 319
rect 1926 323 1935 327
rect 1925 315 1935 319
rect 1789 251 1798 255
rect 3054 269 3058 278
rect 3062 268 3066 278
rect 1789 243 1798 247
rect 1926 251 1935 255
rect 3125 269 3129 278
rect 3133 269 3137 278
rect 3161 269 3165 278
rect 3169 268 3173 278
rect 1926 243 1935 247
rect 3233 269 3237 278
rect 3241 269 3245 278
rect 3269 269 3273 278
rect 3277 268 3281 278
rect 3305 268 3309 278
rect 3313 269 3317 278
rect 3321 268 3325 278
rect 3329 269 3333 278
rect 1789 215 1798 219
rect 1926 215 1935 219
rect 1789 207 1799 211
rect 1925 207 1935 211
rect 1789 179 1799 183
rect 1925 179 1935 183
rect 1789 171 1798 175
rect 1926 171 1935 175
rect 1789 161 1799 165
rect 1925 161 1935 165
rect 1789 153 1798 157
rect 1926 153 1935 157
rect 1789 145 1799 149
rect 1925 145 1935 149
rect 1278 74 1282 83
rect 1286 73 1290 83
rect 1789 137 1798 141
rect 1926 137 1935 141
rect 1349 74 1353 83
rect 1357 74 1361 83
rect 1385 74 1389 83
rect 1393 73 1397 83
rect 3054 127 3058 136
rect 3062 127 3066 137
rect 3125 127 3129 136
rect 3133 127 3137 136
rect 3161 127 3165 136
rect 3169 127 3173 137
rect 1457 74 1461 83
rect 1465 74 1469 83
rect 1493 74 1497 83
rect 1501 73 1505 83
rect 1529 73 1533 83
rect 1537 74 1541 83
rect 1547 73 1551 83
rect 1555 74 1559 83
rect 1563 73 1567 83
rect 1571 74 1575 83
rect 3233 127 3237 136
rect 3241 127 3245 136
rect 3269 127 3273 136
rect 3277 127 3281 137
rect 3305 127 3309 137
rect 3313 127 3317 136
rect 3324 127 3328 137
rect 3332 127 3336 136
rect 1278 -50 1282 -41
rect 1286 -50 1290 -40
rect 1349 -50 1353 -41
rect 1357 -50 1361 -41
rect 1385 -50 1389 -41
rect 1393 -50 1397 -40
rect 1457 -50 1461 -41
rect 1465 -50 1469 -41
rect 1493 -50 1497 -41
rect 1501 -50 1505 -40
rect 1529 -50 1533 -40
rect 1537 -50 1541 -41
rect 1547 -50 1551 -40
rect 1555 -50 1559 -41
rect 1563 -50 1567 -40
rect 1571 -50 1575 -41
rect 1747 -39 1757 -35
rect 1747 -47 1757 -43
rect 1835 -39 1845 -35
rect 1835 -47 1845 -43
rect 1924 -39 1934 -35
rect 1924 -47 1934 -43
rect 2012 -39 2022 -35
rect 2262 -35 2267 -31
rect 2012 -47 2022 -43
rect 2458 -51 2462 -41
rect 2466 -51 2470 -41
rect 2536 -42 2540 -32
rect 2544 -42 2548 -34
rect 2552 -42 2556 -32
rect 2560 -42 2564 -34
rect 2277 -55 2282 -51
rect 2252 -65 2257 -61
rect 2057 -96 2062 -92
rect 2277 -97 2282 -93
rect 1738 -117 1748 -113
rect 1826 -117 1836 -113
rect 1915 -117 1925 -113
rect 2003 -117 2013 -113
rect 2042 -116 2047 -112
rect 2252 -113 2257 -109
rect 2318 -113 2323 -109
rect 1740 -125 1748 -121
rect 1828 -125 1836 -121
rect 1917 -125 1925 -121
rect 2005 -125 2013 -121
rect 2057 -125 2062 -121
rect 2155 -125 2160 -121
rect 1738 -133 1748 -129
rect 1826 -133 1836 -129
rect 1915 -133 1925 -129
rect 2003 -133 2013 -129
rect 1740 -141 1748 -137
rect 1828 -141 1836 -137
rect 1917 -141 1925 -137
rect 2005 -141 2013 -137
rect 2042 -145 2047 -141
rect 2140 -145 2145 -141
rect 2277 -145 2282 -141
rect 2293 -145 2298 -141
rect 3053 -154 3057 -145
rect 3061 -154 3065 -144
rect 3124 -154 3128 -145
rect 3132 -154 3136 -145
rect 3160 -154 3164 -145
rect 3168 -154 3172 -144
rect 3232 -154 3236 -145
rect 3240 -154 3244 -145
rect 3268 -154 3272 -145
rect 3276 -154 3280 -144
rect 3304 -154 3308 -144
rect 3312 -154 3316 -145
rect 3321 -154 3325 -144
rect 3329 -154 3333 -145
rect 2458 -237 2462 -227
rect 2466 -237 2470 -227
rect 2536 -228 2540 -218
rect 2544 -228 2548 -220
rect 2552 -228 2556 -218
rect 2560 -228 2564 -220
rect 1273 -347 1277 -338
rect 1281 -348 1285 -338
rect 1344 -347 1348 -338
rect 1352 -347 1356 -338
rect 1380 -347 1384 -338
rect 1388 -348 1392 -338
rect 1718 -310 1722 -305
rect 1774 -310 1778 -305
rect 1742 -321 1746 -315
rect 1827 -310 1831 -305
rect 1798 -321 1802 -315
rect 1883 -310 1887 -305
rect 1850 -321 1854 -315
rect 1906 -321 1910 -315
rect 1926 -321 1930 -315
rect 2066 -313 2071 -309
rect 1944 -321 1948 -315
rect 1452 -347 1456 -338
rect 1460 -347 1464 -338
rect 1488 -347 1492 -338
rect 1496 -348 1500 -338
rect 1524 -348 1528 -338
rect 1532 -347 1536 -338
rect 1542 -348 1546 -338
rect 1550 -347 1554 -338
rect 1558 -348 1562 -338
rect 1566 -347 1570 -338
rect 2031 -357 2036 -353
rect 2066 -367 2071 -363
rect 2031 -411 2036 -407
rect 2458 -452 2462 -442
rect 2466 -452 2470 -442
rect 2536 -443 2540 -433
rect 2544 -443 2548 -435
rect 2552 -443 2556 -433
rect 2560 -443 2564 -435
rect 1273 -484 1277 -475
rect 1281 -484 1285 -474
rect 1344 -484 1348 -475
rect 1352 -484 1356 -475
rect 1380 -484 1384 -475
rect 1388 -484 1392 -474
rect 1452 -484 1456 -475
rect 1460 -484 1464 -475
rect 1488 -484 1492 -475
rect 1496 -484 1500 -474
rect 1524 -484 1528 -474
rect 1532 -484 1536 -475
rect 1542 -484 1546 -474
rect 1550 -484 1554 -475
rect 1558 -484 1562 -474
rect 1566 -484 1570 -475
rect 3054 -477 3058 -468
rect 3062 -478 3066 -468
rect 3125 -477 3129 -468
rect 3133 -477 3137 -468
rect 3161 -477 3165 -468
rect 3169 -478 3173 -468
rect 3233 -477 3237 -468
rect 3241 -477 3245 -468
rect 3269 -477 3273 -468
rect 3277 -478 3281 -468
rect 3305 -478 3309 -468
rect 3313 -477 3317 -468
rect 3321 -478 3325 -468
rect 3329 -477 3333 -468
rect 1767 -515 1776 -511
rect 1904 -515 1913 -511
rect 1767 -523 1777 -519
rect 1903 -523 1913 -519
rect 1767 -531 1776 -527
rect 1904 -531 1913 -527
rect 1767 -539 1777 -535
rect 1903 -539 1913 -535
rect 1767 -549 1776 -545
rect 1904 -549 1913 -545
rect 1767 -557 1777 -553
rect 1903 -557 1913 -553
rect 1767 -585 1777 -581
rect 1903 -585 1913 -581
rect 1767 -593 1776 -589
rect 1904 -593 1913 -589
rect 1767 -621 1776 -617
rect 1767 -629 1776 -625
rect 1904 -621 1913 -617
rect 1904 -629 1913 -625
rect 3054 -619 3058 -610
rect 3062 -619 3066 -609
rect 3125 -619 3129 -610
rect 3133 -619 3137 -610
rect 3161 -619 3165 -610
rect 3169 -619 3173 -609
rect 3233 -619 3237 -610
rect 3241 -619 3245 -610
rect 3269 -619 3273 -610
rect 3277 -619 3281 -609
rect 3305 -619 3309 -609
rect 3313 -619 3317 -610
rect 3321 -619 3325 -609
rect 3329 -619 3333 -610
rect 1767 -693 1777 -689
rect 1767 -701 1776 -697
rect 1903 -693 1913 -689
rect 1904 -701 1913 -697
rect 1767 -729 1776 -725
rect 1904 -729 1913 -725
rect 1767 -737 1776 -733
rect 1904 -737 1913 -733
rect 1767 -800 1777 -796
rect 1767 -808 1776 -804
rect 1903 -800 1913 -796
rect 1904 -808 1913 -804
<< pdcontact >>
rect 1756 503 1776 507
rect 1948 503 1968 507
rect 1756 495 1776 499
rect 1948 495 1968 499
rect 1756 467 1776 471
rect 1948 467 1968 471
rect 1756 459 1776 463
rect 1948 459 1968 463
rect 1756 395 1776 399
rect 1756 387 1776 391
rect 1948 395 1968 399
rect 1948 387 1968 391
rect 1756 287 1776 291
rect 1948 287 1968 291
rect 2981 291 2985 311
rect 2989 291 2993 311
rect 3017 291 3021 311
rect 3025 291 3029 311
rect 1756 279 1776 283
rect 1948 279 1968 283
rect 3089 291 3093 311
rect 3097 291 3101 311
rect 3197 291 3201 311
rect 3205 291 3209 311
rect 3305 291 3309 311
rect 3313 291 3317 311
rect 3321 291 3325 311
rect 3329 291 3333 311
rect 1756 179 1776 183
rect 1948 179 1968 183
rect 1756 171 1776 175
rect 1948 171 1968 175
rect 1756 161 1776 165
rect 1948 161 1968 165
rect 1756 153 1776 157
rect 1948 153 1968 157
rect 1756 145 1776 149
rect 1948 145 1968 149
rect 1205 96 1209 116
rect 1213 96 1217 116
rect 1241 96 1245 116
rect 1249 96 1253 116
rect 1313 96 1317 116
rect 1321 96 1325 116
rect 1756 137 1776 141
rect 1948 137 1968 141
rect 1421 96 1425 116
rect 1429 96 1433 116
rect 1529 96 1533 116
rect 1537 96 1541 116
rect 1547 96 1551 116
rect 1555 96 1559 116
rect 1563 96 1567 116
rect 1571 96 1575 116
rect 2981 94 2985 114
rect 2989 94 2993 114
rect 3017 94 3021 114
rect 3025 94 3029 114
rect 3089 94 3093 114
rect 3097 94 3101 114
rect 3197 94 3201 114
rect 3205 94 3209 114
rect 3305 94 3309 114
rect 3313 94 3317 114
rect 3324 94 3328 114
rect 3332 94 3336 114
rect 2467 -5 2517 -1
rect 2467 -13 2517 -9
rect 2536 -17 2540 3
rect 2544 -17 2548 3
rect 2552 -17 2556 3
rect 2560 -17 2564 3
rect 1205 -83 1209 -63
rect 1213 -83 1217 -63
rect 1241 -83 1245 -63
rect 1249 -83 1253 -63
rect 1313 -83 1317 -63
rect 1321 -83 1325 -63
rect 2467 -21 2517 -17
rect 2467 -29 2517 -25
rect 1421 -83 1425 -63
rect 1429 -83 1433 -63
rect 1529 -83 1533 -63
rect 1537 -83 1541 -63
rect 1547 -83 1551 -63
rect 1555 -83 1559 -63
rect 1563 -83 1567 -63
rect 1571 -83 1575 -63
rect 1707 -94 1711 -44
rect 1715 -94 1719 -44
rect 1723 -94 1727 -44
rect 1731 -94 1735 -44
rect 1795 -94 1799 -44
rect 1803 -94 1807 -44
rect 1811 -94 1815 -44
rect 1819 -94 1823 -44
rect 2208 -35 2214 -31
rect 1884 -94 1888 -44
rect 1892 -94 1896 -44
rect 1900 -94 1904 -44
rect 1908 -94 1912 -44
rect 1972 -94 1976 -44
rect 1980 -94 1984 -44
rect 1988 -94 1992 -44
rect 1996 -94 2000 -44
rect 2222 -45 2228 -41
rect 2208 -55 2214 -51
rect 2222 -65 2228 -61
rect 2208 -75 2214 -71
rect 2222 -87 2228 -83
rect 2111 -96 2117 -92
rect 2208 -97 2214 -93
rect 2097 -106 2103 -102
rect 1703 -117 1723 -113
rect 1791 -117 1811 -113
rect 1880 -117 1900 -113
rect 1968 -117 1988 -113
rect 2111 -116 2117 -112
rect 2222 -113 2228 -109
rect 2346 -113 2352 -109
rect 1703 -125 1723 -121
rect 1791 -125 1811 -121
rect 1880 -125 1900 -121
rect 1968 -125 1988 -121
rect 2111 -125 2117 -121
rect 2192 -125 2198 -121
rect 2208 -123 2214 -119
rect 2360 -123 2366 -119
rect 1703 -133 1723 -129
rect 1791 -133 1811 -129
rect 1880 -133 1900 -129
rect 1968 -133 1988 -129
rect 1703 -141 1723 -137
rect 1791 -141 1811 -137
rect 1880 -141 1900 -137
rect 1968 -141 1988 -137
rect 2097 -135 2103 -131
rect 2178 -135 2184 -131
rect 2222 -135 2228 -131
rect 2346 -135 2352 -131
rect 2111 -145 2117 -141
rect 2192 -145 2198 -141
rect 2208 -145 2214 -141
rect 2360 -145 2366 -141
rect 2467 -191 2517 -187
rect 2467 -199 2517 -195
rect 2536 -203 2540 -183
rect 2544 -203 2548 -183
rect 2552 -203 2556 -183
rect 2560 -203 2564 -183
rect 2980 -187 2984 -167
rect 2988 -187 2992 -167
rect 3016 -187 3020 -167
rect 3024 -187 3028 -167
rect 3088 -187 3092 -167
rect 3096 -187 3100 -167
rect 3196 -187 3200 -167
rect 3204 -187 3208 -167
rect 2467 -207 2517 -203
rect 3304 -187 3308 -167
rect 3312 -187 3316 -167
rect 3321 -187 3325 -167
rect 3329 -187 3333 -167
rect 2467 -215 2517 -211
rect 1200 -325 1204 -305
rect 1208 -325 1212 -305
rect 1236 -325 1240 -305
rect 1244 -325 1248 -305
rect 1308 -325 1312 -305
rect 1316 -325 1320 -305
rect 1416 -325 1420 -305
rect 1424 -325 1428 -305
rect 1524 -325 1528 -305
rect 1532 -325 1536 -305
rect 1542 -325 1546 -305
rect 1550 -325 1554 -305
rect 1558 -325 1562 -305
rect 1566 -325 1570 -305
rect 1973 -313 1979 -309
rect 1987 -323 1993 -319
rect 1973 -335 1979 -331
rect 1698 -356 1702 -350
rect 1708 -342 1712 -336
rect 1718 -356 1722 -350
rect 1734 -356 1738 -350
rect 1742 -342 1746 -336
rect 1754 -356 1758 -350
rect 1764 -342 1768 -336
rect 1774 -356 1778 -350
rect 1790 -356 1794 -350
rect 1798 -342 1802 -336
rect 1807 -356 1811 -350
rect 1817 -342 1821 -336
rect 1827 -356 1831 -350
rect 1842 -356 1846 -350
rect 1850 -342 1854 -336
rect 1863 -356 1867 -350
rect 1873 -342 1877 -336
rect 1883 -356 1887 -350
rect 1898 -356 1902 -350
rect 1906 -342 1910 -336
rect 1918 -356 1922 -350
rect 1926 -342 1930 -336
rect 1936 -356 1940 -350
rect 1944 -342 1948 -336
rect 1987 -347 1993 -343
rect 1973 -357 1979 -353
rect 1973 -367 1979 -363
rect 1987 -377 1993 -373
rect 1973 -389 1979 -385
rect 1987 -401 1993 -397
rect 1973 -411 1979 -407
rect 2467 -406 2517 -402
rect 2467 -414 2517 -410
rect 2536 -418 2540 -398
rect 2544 -418 2548 -398
rect 2552 -418 2556 -398
rect 2560 -418 2564 -398
rect 2467 -422 2517 -418
rect 2467 -430 2517 -426
rect 1200 -517 1204 -497
rect 1208 -517 1212 -497
rect 1236 -517 1240 -497
rect 1244 -517 1248 -497
rect 1308 -517 1312 -497
rect 1316 -517 1320 -497
rect 2981 -455 2985 -435
rect 2989 -455 2993 -435
rect 3017 -455 3021 -435
rect 3025 -455 3029 -435
rect 1416 -517 1420 -497
rect 1424 -517 1428 -497
rect 3089 -455 3093 -435
rect 3097 -455 3101 -435
rect 1524 -517 1528 -497
rect 1532 -517 1536 -497
rect 1542 -517 1546 -497
rect 1550 -517 1554 -497
rect 1558 -517 1562 -497
rect 1566 -517 1570 -497
rect 3197 -455 3201 -435
rect 3205 -455 3209 -435
rect 3305 -455 3309 -435
rect 3313 -455 3317 -435
rect 3321 -455 3325 -435
rect 3329 -455 3333 -435
rect 1734 -515 1754 -511
rect 1926 -515 1946 -511
rect 1734 -523 1754 -519
rect 1926 -523 1946 -519
rect 1734 -531 1754 -527
rect 1926 -531 1946 -527
rect 1734 -539 1754 -535
rect 1926 -539 1946 -535
rect 1734 -549 1754 -545
rect 1926 -549 1946 -545
rect 1734 -557 1754 -553
rect 1926 -557 1946 -553
rect 2981 -652 2985 -632
rect 2989 -652 2993 -632
rect 3017 -652 3021 -632
rect 3025 -652 3029 -632
rect 1734 -657 1754 -653
rect 1926 -657 1946 -653
rect 3089 -652 3093 -632
rect 3097 -652 3101 -632
rect 1734 -665 1754 -661
rect 1926 -665 1946 -661
rect 3197 -652 3201 -632
rect 3205 -652 3209 -632
rect 3305 -652 3309 -632
rect 3313 -652 3317 -632
rect 3321 -652 3325 -632
rect 3329 -652 3333 -632
rect 1734 -765 1754 -761
rect 1734 -773 1754 -769
rect 1926 -765 1946 -761
rect 1926 -773 1946 -769
rect 1734 -837 1754 -833
rect 1926 -837 1946 -833
rect 1734 -845 1754 -841
rect 1926 -845 1946 -841
rect 1734 -873 1754 -869
rect 1926 -873 1946 -869
rect 1734 -881 1754 -877
rect 1926 -881 1946 -877
<< psubstratepdiff >>
rect 3317 260 3320 264
rect 1803 166 1807 167
rect 1917 166 1921 167
rect 3321 141 3323 145
rect 1545 65 1546 69
rect 1545 -36 1546 -32
rect 1540 -356 1541 -352
rect 1540 -470 1541 -466
rect 1781 -541 1785 -540
rect 1895 -541 1899 -540
<< nsubstratendiff >>
rect 3322 86 3323 90
<< psubstratepcontact >>
rect 1803 513 1807 517
rect 1917 513 1921 517
rect 1803 504 1807 508
rect 1917 504 1921 508
rect 1803 487 1807 491
rect 1917 487 1921 491
rect 1803 477 1807 481
rect 1917 477 1921 481
rect 1803 468 1807 472
rect 1917 468 1921 472
rect 1803 451 1807 455
rect 1917 451 1921 455
rect 1803 441 1807 445
rect 1917 441 1921 445
rect 1803 432 1807 436
rect 1917 432 1921 436
rect 1803 415 1807 419
rect 1917 415 1921 419
rect 1803 405 1807 409
rect 1917 405 1921 409
rect 1803 396 1807 400
rect 1917 396 1921 400
rect 1803 379 1807 383
rect 1917 379 1921 383
rect 1803 369 1807 373
rect 1917 369 1921 373
rect 1803 360 1807 364
rect 1917 360 1921 364
rect 1803 343 1807 347
rect 1917 343 1921 347
rect 1803 333 1807 337
rect 1917 333 1921 337
rect 1803 324 1807 328
rect 1917 324 1921 328
rect 1803 307 1807 311
rect 1917 307 1921 311
rect 1803 297 1807 301
rect 1917 297 1921 301
rect 1803 288 1807 292
rect 1917 288 1921 292
rect 1803 271 1807 275
rect 1917 271 1921 275
rect 1803 261 1807 265
rect 1917 261 1921 265
rect 2971 260 2975 264
rect 2980 260 2984 264
rect 1803 252 1807 256
rect 1917 252 1921 256
rect 2997 260 3001 264
rect 3007 260 3011 264
rect 3016 260 3020 264
rect 3033 260 3037 264
rect 3043 260 3047 264
rect 3052 260 3056 264
rect 3069 260 3073 264
rect 3079 260 3083 264
rect 3088 260 3092 264
rect 3105 260 3109 264
rect 3115 260 3119 264
rect 3124 260 3128 264
rect 3141 260 3145 264
rect 3151 260 3155 264
rect 3160 260 3164 264
rect 3177 260 3181 264
rect 3187 260 3191 264
rect 3196 260 3200 264
rect 3213 260 3217 264
rect 3223 260 3227 264
rect 3232 260 3236 264
rect 3249 260 3253 264
rect 3259 260 3263 264
rect 3268 260 3272 264
rect 3285 260 3289 264
rect 3295 260 3299 264
rect 3304 260 3308 264
rect 3320 260 3324 264
rect 1803 235 1807 239
rect 1917 235 1921 239
rect 1803 225 1807 229
rect 1917 225 1921 229
rect 1803 216 1807 220
rect 1917 216 1921 220
rect 1803 199 1807 203
rect 1917 199 1921 203
rect 1803 189 1807 193
rect 1917 189 1921 193
rect 1803 180 1807 184
rect 1917 180 1921 184
rect 1803 162 1807 166
rect 1917 162 1921 166
rect 1803 146 1807 150
rect 1917 146 1921 150
rect 1195 65 1199 69
rect 1204 65 1208 69
rect 1221 65 1225 69
rect 1231 65 1235 69
rect 1240 65 1244 69
rect 1257 65 1261 69
rect 1267 65 1271 69
rect 1276 65 1280 69
rect 1293 65 1297 69
rect 1303 65 1307 69
rect 1312 65 1316 69
rect 2971 141 2975 145
rect 2980 141 2984 145
rect 1329 65 1333 69
rect 1339 65 1343 69
rect 1348 65 1352 69
rect 1365 65 1369 69
rect 1375 65 1379 69
rect 1384 65 1388 69
rect 1401 65 1405 69
rect 1411 65 1415 69
rect 1420 65 1424 69
rect 1803 129 1807 133
rect 1917 129 1921 133
rect 2997 141 3001 145
rect 3007 141 3011 145
rect 3016 141 3020 145
rect 3033 141 3037 145
rect 3043 141 3047 145
rect 3052 141 3056 145
rect 3069 141 3073 145
rect 3079 141 3083 145
rect 3088 141 3092 145
rect 3105 141 3109 145
rect 3115 141 3119 145
rect 3124 141 3128 145
rect 3141 141 3145 145
rect 3151 141 3155 145
rect 3160 141 3164 145
rect 3177 141 3181 145
rect 3187 141 3191 145
rect 3196 141 3200 145
rect 3213 141 3217 145
rect 3223 141 3227 145
rect 3232 141 3236 145
rect 3249 141 3253 145
rect 3259 141 3263 145
rect 3268 141 3272 145
rect 3285 141 3289 145
rect 3295 141 3299 145
rect 3304 141 3308 145
rect 3323 141 3327 145
rect 3340 141 3344 145
rect 1437 65 1441 69
rect 1447 65 1451 69
rect 1456 65 1460 69
rect 1473 65 1477 69
rect 1483 65 1487 69
rect 1492 65 1496 69
rect 1509 65 1513 69
rect 1519 65 1523 69
rect 1528 65 1532 69
rect 1546 65 1550 69
rect 1562 65 1566 69
rect 1579 65 1583 69
rect 1195 -36 1199 -32
rect 1204 -36 1208 -32
rect 1221 -36 1225 -32
rect 1231 -36 1235 -32
rect 1240 -36 1244 -32
rect 1257 -36 1261 -32
rect 1267 -36 1271 -32
rect 1276 -36 1280 -32
rect 1293 -36 1297 -32
rect 1303 -36 1307 -32
rect 1312 -36 1316 -32
rect 1329 -36 1333 -32
rect 1339 -36 1343 -32
rect 1348 -36 1352 -32
rect 1365 -36 1369 -32
rect 1375 -36 1379 -32
rect 1384 -36 1388 -32
rect 1401 -36 1405 -32
rect 1411 -36 1415 -32
rect 1420 -36 1424 -32
rect 1437 -36 1441 -32
rect 1447 -36 1451 -32
rect 1456 -36 1460 -32
rect 1473 -36 1477 -32
rect 1483 -36 1487 -32
rect 1492 -36 1496 -32
rect 1509 -36 1513 -32
rect 1519 -36 1523 -32
rect 1528 -36 1532 -32
rect 1546 -36 1550 -32
rect 1562 -36 1566 -32
rect 1579 -36 1583 -32
rect 2970 -140 2974 -136
rect 2979 -140 2983 -136
rect 2996 -140 3000 -136
rect 3006 -140 3010 -136
rect 3015 -140 3019 -136
rect 3032 -140 3036 -136
rect 3042 -140 3046 -136
rect 3051 -140 3055 -136
rect 3068 -140 3072 -136
rect 3078 -140 3082 -136
rect 3087 -140 3091 -136
rect 3104 -140 3108 -136
rect 3114 -140 3118 -136
rect 3123 -140 3127 -136
rect 3140 -140 3144 -136
rect 3150 -140 3154 -136
rect 3159 -140 3163 -136
rect 3176 -140 3180 -136
rect 3186 -140 3190 -136
rect 3195 -140 3199 -136
rect 3212 -140 3216 -136
rect 3222 -140 3226 -136
rect 3231 -140 3235 -136
rect 3248 -140 3252 -136
rect 3258 -140 3262 -136
rect 3267 -140 3271 -136
rect 3284 -140 3288 -136
rect 3294 -140 3298 -136
rect 3303 -140 3307 -136
rect 3320 -140 3324 -136
rect 3337 -140 3341 -136
rect 1190 -356 1194 -352
rect 1199 -356 1203 -352
rect 1216 -356 1220 -352
rect 1226 -356 1230 -352
rect 1235 -356 1239 -352
rect 1252 -356 1256 -352
rect 1262 -356 1266 -352
rect 1271 -356 1275 -352
rect 1288 -356 1292 -352
rect 1298 -356 1302 -352
rect 1307 -356 1311 -352
rect 1324 -356 1328 -352
rect 1334 -356 1338 -352
rect 1343 -356 1347 -352
rect 1360 -356 1364 -352
rect 1370 -356 1374 -352
rect 1379 -356 1383 -352
rect 1396 -356 1400 -352
rect 1406 -356 1410 -352
rect 1415 -356 1419 -352
rect 1432 -356 1436 -352
rect 1442 -356 1446 -352
rect 1451 -356 1455 -352
rect 1468 -356 1472 -352
rect 1478 -356 1482 -352
rect 1487 -356 1491 -352
rect 1504 -356 1508 -352
rect 1514 -356 1518 -352
rect 1523 -356 1527 -352
rect 1541 -356 1545 -352
rect 1557 -356 1561 -352
rect 1574 -356 1578 -352
rect 1190 -470 1194 -466
rect 1199 -470 1203 -466
rect 1216 -470 1220 -466
rect 1226 -470 1230 -466
rect 1235 -470 1239 -466
rect 1252 -470 1256 -466
rect 1262 -470 1266 -466
rect 1271 -470 1275 -466
rect 1288 -470 1292 -466
rect 1298 -470 1302 -466
rect 1307 -470 1311 -466
rect 1324 -470 1328 -466
rect 1334 -470 1338 -466
rect 1343 -470 1347 -466
rect 1360 -470 1364 -466
rect 1370 -470 1374 -466
rect 1379 -470 1383 -466
rect 1396 -470 1400 -466
rect 1406 -470 1410 -466
rect 1415 -470 1419 -466
rect 1432 -470 1436 -466
rect 1442 -470 1446 -466
rect 1451 -470 1455 -466
rect 1468 -470 1472 -466
rect 1478 -470 1482 -466
rect 1487 -470 1491 -466
rect 1504 -470 1508 -466
rect 1514 -470 1518 -466
rect 1523 -470 1527 -466
rect 1541 -470 1545 -466
rect 1557 -470 1561 -466
rect 1574 -470 1578 -466
rect 2971 -486 2975 -482
rect 2980 -486 2984 -482
rect 2997 -486 3001 -482
rect 3007 -486 3011 -482
rect 3016 -486 3020 -482
rect 3033 -486 3037 -482
rect 3043 -486 3047 -482
rect 3052 -486 3056 -482
rect 3069 -486 3073 -482
rect 3079 -486 3083 -482
rect 3088 -486 3092 -482
rect 3105 -486 3109 -482
rect 3115 -486 3119 -482
rect 3124 -486 3128 -482
rect 3141 -486 3145 -482
rect 3151 -486 3155 -482
rect 3160 -486 3164 -482
rect 3177 -486 3181 -482
rect 3187 -486 3191 -482
rect 3196 -486 3200 -482
rect 3213 -486 3217 -482
rect 3223 -486 3227 -482
rect 3232 -486 3236 -482
rect 3249 -486 3253 -482
rect 3259 -486 3263 -482
rect 3268 -486 3272 -482
rect 3285 -486 3289 -482
rect 3295 -486 3299 -482
rect 3304 -486 3308 -482
rect 3320 -486 3324 -482
rect 3337 -486 3341 -482
rect 1781 -507 1785 -503
rect 1895 -507 1899 -503
rect 1781 -524 1785 -520
rect 1895 -524 1899 -520
rect 1781 -540 1785 -536
rect 1895 -540 1899 -536
rect 1781 -558 1785 -554
rect 1895 -558 1899 -554
rect 1781 -567 1785 -563
rect 1895 -567 1899 -563
rect 1781 -577 1785 -573
rect 1895 -577 1899 -573
rect 1781 -594 1785 -590
rect 1895 -594 1899 -590
rect 1781 -603 1785 -599
rect 1895 -603 1899 -599
rect 2971 -605 2975 -601
rect 2980 -605 2984 -601
rect 1781 -613 1785 -609
rect 1895 -613 1899 -609
rect 1781 -630 1785 -626
rect 1895 -630 1899 -626
rect 2997 -605 3001 -601
rect 3007 -605 3011 -601
rect 3016 -605 3020 -601
rect 3033 -605 3037 -601
rect 3043 -605 3047 -601
rect 3052 -605 3056 -601
rect 3069 -605 3073 -601
rect 3079 -605 3083 -601
rect 3088 -605 3092 -601
rect 1781 -639 1785 -635
rect 1895 -639 1899 -635
rect 1781 -649 1785 -645
rect 1895 -649 1899 -645
rect 3105 -605 3109 -601
rect 3115 -605 3119 -601
rect 3124 -605 3128 -601
rect 3141 -605 3145 -601
rect 3151 -605 3155 -601
rect 3160 -605 3164 -601
rect 3177 -605 3181 -601
rect 3187 -605 3191 -601
rect 3196 -605 3200 -601
rect 1781 -666 1785 -662
rect 1895 -666 1899 -662
rect 3213 -605 3217 -601
rect 3223 -605 3227 -601
rect 3232 -605 3236 -601
rect 3249 -605 3253 -601
rect 3259 -605 3263 -601
rect 3268 -605 3272 -601
rect 3285 -605 3289 -601
rect 3295 -605 3299 -601
rect 3304 -605 3308 -601
rect 3320 -605 3324 -601
rect 3337 -605 3341 -601
rect 1781 -675 1785 -671
rect 1895 -675 1899 -671
rect 1781 -685 1785 -681
rect 1895 -685 1899 -681
rect 1781 -702 1785 -698
rect 1895 -702 1899 -698
rect 1781 -711 1785 -707
rect 1895 -711 1899 -707
rect 1781 -721 1785 -717
rect 1895 -721 1899 -717
rect 1781 -738 1785 -734
rect 1895 -738 1899 -734
rect 1781 -747 1785 -743
rect 1895 -747 1899 -743
rect 1781 -757 1785 -753
rect 1895 -757 1899 -753
rect 1781 -774 1785 -770
rect 1895 -774 1899 -770
rect 1781 -783 1785 -779
rect 1895 -783 1899 -779
rect 1781 -793 1785 -789
rect 1895 -793 1899 -789
rect 1781 -810 1785 -806
rect 1895 -810 1899 -806
rect 1781 -819 1785 -815
rect 1895 -819 1899 -815
rect 1781 -829 1785 -825
rect 1895 -829 1899 -825
rect 1781 -846 1785 -842
rect 1895 -846 1899 -842
rect 1781 -855 1785 -851
rect 1895 -855 1899 -851
rect 1781 -865 1785 -861
rect 1895 -865 1899 -861
rect 1781 -882 1785 -878
rect 1895 -882 1899 -878
rect 1781 -891 1785 -887
rect 1895 -891 1899 -887
<< nsubstratencontact >>
rect 1748 512 1752 516
rect 1972 512 1976 516
rect 1748 504 1752 508
rect 1972 504 1976 508
rect 1748 495 1752 499
rect 1972 495 1976 499
rect 1748 486 1752 490
rect 1972 486 1976 490
rect 1748 476 1752 480
rect 1972 476 1976 480
rect 1748 468 1752 472
rect 1972 468 1976 472
rect 1748 459 1752 463
rect 1972 459 1976 463
rect 1748 450 1752 454
rect 1972 450 1976 454
rect 1748 423 1752 427
rect 1972 423 1976 427
rect 1748 414 1752 418
rect 1972 414 1976 418
rect 1748 404 1752 408
rect 1972 404 1976 408
rect 1748 396 1752 400
rect 1748 387 1752 391
rect 1972 396 1976 400
rect 1972 387 1976 391
rect 1748 378 1752 382
rect 1972 378 1976 382
rect 1748 368 1752 372
rect 1972 368 1976 372
rect 1748 360 1752 364
rect 1972 360 1976 364
rect 1748 351 1752 355
rect 1972 351 1976 355
rect 1748 342 1752 346
rect 1972 342 1976 346
rect 1748 315 1752 319
rect 1972 315 1976 319
rect 2972 315 2976 319
rect 2980 315 2984 319
rect 2989 315 2993 319
rect 2998 315 3002 319
rect 3008 315 3012 319
rect 3016 315 3020 319
rect 3025 315 3029 319
rect 3034 315 3038 319
rect 3061 315 3065 319
rect 3070 315 3074 319
rect 3080 315 3084 319
rect 3088 315 3092 319
rect 3097 315 3101 319
rect 3106 315 3110 319
rect 3116 315 3120 319
rect 3124 315 3128 319
rect 1748 306 1752 310
rect 1972 306 1976 310
rect 1748 296 1752 300
rect 1972 296 1976 300
rect 1748 288 1752 292
rect 1972 288 1976 292
rect 1748 279 1752 283
rect 1972 279 1976 283
rect 1748 270 1752 274
rect 1972 270 1976 274
rect 1748 243 1752 247
rect 3133 315 3137 319
rect 3142 315 3146 319
rect 3169 315 3173 319
rect 3178 315 3182 319
rect 3188 315 3192 319
rect 3196 315 3200 319
rect 3205 315 3209 319
rect 3214 315 3218 319
rect 3241 315 3245 319
rect 3250 315 3254 319
rect 3260 315 3264 319
rect 3268 315 3272 319
rect 1972 243 1976 247
rect 3277 315 3281 319
rect 3286 315 3290 319
rect 3296 315 3300 319
rect 3304 315 3308 319
rect 3329 315 3333 319
rect 1748 234 1752 238
rect 1972 234 1976 238
rect 1748 224 1752 228
rect 1972 224 1976 228
rect 1748 216 1752 220
rect 1972 216 1976 220
rect 1748 207 1752 211
rect 1972 207 1976 211
rect 1748 198 1752 202
rect 1972 198 1976 202
rect 1748 188 1752 192
rect 1972 188 1976 192
rect 1748 180 1752 184
rect 1972 180 1976 184
rect 1748 171 1752 175
rect 1972 171 1976 175
rect 1748 162 1752 166
rect 1972 162 1976 166
rect 1748 153 1752 157
rect 1972 153 1976 157
rect 1196 120 1200 124
rect 1204 120 1208 124
rect 1213 120 1217 124
rect 1222 120 1226 124
rect 1232 120 1236 124
rect 1240 120 1244 124
rect 1249 120 1253 124
rect 1258 120 1262 124
rect 1285 120 1289 124
rect 1294 120 1298 124
rect 1304 120 1308 124
rect 1312 120 1316 124
rect 1321 120 1325 124
rect 1330 120 1334 124
rect 1340 120 1344 124
rect 1348 120 1352 124
rect 1357 120 1361 124
rect 1366 120 1370 124
rect 1393 120 1397 124
rect 1402 120 1406 124
rect 1412 120 1416 124
rect 1420 120 1424 124
rect 1748 137 1752 141
rect 1972 137 1976 141
rect 1429 120 1433 124
rect 1438 120 1442 124
rect 1465 120 1469 124
rect 1474 120 1478 124
rect 1484 120 1488 124
rect 1492 120 1496 124
rect 1501 120 1505 124
rect 1510 120 1514 124
rect 1520 120 1524 124
rect 1528 120 1532 124
rect 1748 128 1752 132
rect 1972 128 1976 132
rect 1537 120 1541 124
rect 1546 120 1550 124
rect 1555 120 1559 124
rect 1571 120 1575 124
rect 1580 120 1584 124
rect 2972 86 2976 90
rect 2980 86 2984 90
rect 2989 86 2993 90
rect 2998 86 3002 90
rect 3008 86 3012 90
rect 3016 86 3020 90
rect 3025 86 3029 90
rect 3034 86 3038 90
rect 3061 86 3065 90
rect 3070 86 3074 90
rect 3080 86 3084 90
rect 3088 86 3092 90
rect 3097 86 3101 90
rect 3106 86 3110 90
rect 3116 86 3120 90
rect 3124 86 3128 90
rect 3133 86 3137 90
rect 3142 86 3146 90
rect 3169 86 3173 90
rect 3178 86 3182 90
rect 3188 86 3192 90
rect 3196 86 3200 90
rect 3205 86 3209 90
rect 3214 86 3218 90
rect 3241 86 3245 90
rect 3250 86 3254 90
rect 3260 86 3264 90
rect 3268 86 3272 90
rect 3277 86 3281 90
rect 3286 86 3290 90
rect 3296 86 3300 90
rect 3304 86 3308 90
rect 3313 86 3317 90
rect 3323 86 3327 90
rect 3332 86 3336 90
rect 3341 86 3345 90
rect 2532 8 2536 12
rect 2545 8 2549 12
rect 2561 8 2565 12
rect 1196 -91 1200 -87
rect 1204 -91 1208 -87
rect 1213 -91 1217 -87
rect 1222 -91 1226 -87
rect 1232 -91 1236 -87
rect 1240 -91 1244 -87
rect 1249 -91 1253 -87
rect 1258 -91 1262 -87
rect 1285 -91 1289 -87
rect 1294 -91 1298 -87
rect 1304 -91 1308 -87
rect 1312 -91 1316 -87
rect 1321 -91 1325 -87
rect 1330 -91 1334 -87
rect 1340 -91 1344 -87
rect 1348 -91 1352 -87
rect 1357 -91 1361 -87
rect 1366 -91 1370 -87
rect 1393 -91 1397 -87
rect 1402 -91 1406 -87
rect 1412 -91 1416 -87
rect 1420 -91 1424 -87
rect 1429 -91 1433 -87
rect 1438 -91 1442 -87
rect 1465 -91 1469 -87
rect 1474 -91 1478 -87
rect 1484 -91 1488 -87
rect 1492 -91 1496 -87
rect 1501 -91 1505 -87
rect 1510 -91 1514 -87
rect 1520 -91 1524 -87
rect 1528 -91 1532 -87
rect 1537 -91 1541 -87
rect 1546 -91 1550 -87
rect 1555 -91 1559 -87
rect 1571 -91 1575 -87
rect 1580 -91 1584 -87
rect 1694 -113 1698 -109
rect 1782 -113 1786 -109
rect 1871 -113 1875 -109
rect 1959 -113 1963 -109
rect 1694 -128 1698 -124
rect 1782 -126 1786 -122
rect 1959 -128 1963 -124
rect 1871 -133 1875 -129
rect 1694 -143 1698 -139
rect 1782 -142 1786 -138
rect 1871 -144 1875 -140
rect 1959 -144 1963 -140
rect 2532 -178 2536 -174
rect 2545 -178 2549 -174
rect 2561 -178 2565 -174
rect 2971 -195 2975 -191
rect 2979 -195 2983 -191
rect 2988 -195 2992 -191
rect 2997 -195 3001 -191
rect 3007 -195 3011 -191
rect 3015 -195 3019 -191
rect 3024 -195 3028 -191
rect 3033 -195 3037 -191
rect 3060 -195 3064 -191
rect 3069 -195 3073 -191
rect 3079 -195 3083 -191
rect 3087 -195 3091 -191
rect 3096 -195 3100 -191
rect 3105 -195 3109 -191
rect 3115 -195 3119 -191
rect 3123 -195 3127 -191
rect 3132 -195 3136 -191
rect 3141 -195 3145 -191
rect 3168 -195 3172 -191
rect 3177 -195 3181 -191
rect 3187 -195 3191 -191
rect 3195 -195 3199 -191
rect 3204 -195 3208 -191
rect 3213 -195 3217 -191
rect 3240 -195 3244 -191
rect 3249 -195 3253 -191
rect 3259 -195 3263 -191
rect 3267 -195 3271 -191
rect 3276 -195 3280 -191
rect 3285 -195 3289 -191
rect 3295 -195 3299 -191
rect 3303 -195 3307 -191
rect 3320 -195 3324 -191
rect 3329 -195 3333 -191
rect 3338 -195 3342 -191
rect 1191 -301 1195 -297
rect 1199 -301 1203 -297
rect 1208 -301 1212 -297
rect 1217 -301 1221 -297
rect 1227 -301 1231 -297
rect 1235 -301 1239 -297
rect 1244 -301 1248 -297
rect 1253 -301 1257 -297
rect 1280 -301 1284 -297
rect 1289 -301 1293 -297
rect 1299 -301 1303 -297
rect 1307 -301 1311 -297
rect 1316 -301 1320 -297
rect 1325 -301 1329 -297
rect 1335 -301 1339 -297
rect 1343 -301 1347 -297
rect 1352 -301 1356 -297
rect 1361 -301 1365 -297
rect 1388 -301 1392 -297
rect 1397 -301 1401 -297
rect 1407 -301 1411 -297
rect 1415 -301 1419 -297
rect 1424 -301 1428 -297
rect 1433 -301 1437 -297
rect 1460 -301 1464 -297
rect 1469 -301 1473 -297
rect 1479 -301 1483 -297
rect 1487 -301 1491 -297
rect 1496 -301 1500 -297
rect 1505 -301 1509 -297
rect 1515 -301 1519 -297
rect 1523 -301 1527 -297
rect 1532 -301 1536 -297
rect 1541 -301 1545 -297
rect 1550 -301 1554 -297
rect 1566 -301 1570 -297
rect 1575 -301 1579 -297
rect 2532 -393 2536 -389
rect 2545 -393 2549 -389
rect 2561 -393 2565 -389
rect 2972 -431 2976 -427
rect 2980 -431 2984 -427
rect 2989 -431 2993 -427
rect 2998 -431 3002 -427
rect 3008 -431 3012 -427
rect 3016 -431 3020 -427
rect 3025 -431 3029 -427
rect 3034 -431 3038 -427
rect 3061 -431 3065 -427
rect 3070 -431 3074 -427
rect 3080 -431 3084 -427
rect 3088 -431 3092 -427
rect 3097 -431 3101 -427
rect 3106 -431 3110 -427
rect 3116 -431 3120 -427
rect 3124 -431 3128 -427
rect 1191 -525 1195 -521
rect 1199 -525 1203 -521
rect 1208 -525 1212 -521
rect 1217 -525 1221 -521
rect 1227 -525 1231 -521
rect 1235 -525 1239 -521
rect 1244 -525 1248 -521
rect 1253 -525 1257 -521
rect 1280 -525 1284 -521
rect 1289 -525 1293 -521
rect 1299 -525 1303 -521
rect 1307 -525 1311 -521
rect 1316 -525 1320 -521
rect 1325 -525 1329 -521
rect 1335 -525 1339 -521
rect 1343 -525 1347 -521
rect 1352 -525 1356 -521
rect 1361 -525 1365 -521
rect 1388 -525 1392 -521
rect 1397 -525 1401 -521
rect 1407 -525 1411 -521
rect 1415 -525 1419 -521
rect 1424 -525 1428 -521
rect 1433 -525 1437 -521
rect 1460 -525 1464 -521
rect 1469 -525 1473 -521
rect 1479 -525 1483 -521
rect 1487 -525 1491 -521
rect 3133 -431 3137 -427
rect 3142 -431 3146 -427
rect 3169 -431 3173 -427
rect 3178 -431 3182 -427
rect 3188 -431 3192 -427
rect 3196 -431 3200 -427
rect 3205 -431 3209 -427
rect 3214 -431 3218 -427
rect 3241 -431 3245 -427
rect 3250 -431 3254 -427
rect 3260 -431 3264 -427
rect 3268 -431 3272 -427
rect 3277 -431 3281 -427
rect 3286 -431 3290 -427
rect 3296 -431 3300 -427
rect 3304 -431 3308 -427
rect 3320 -431 3324 -427
rect 3329 -431 3333 -427
rect 1726 -506 1730 -502
rect 1950 -506 1954 -502
rect 1726 -515 1730 -511
rect 1950 -515 1954 -511
rect 1496 -525 1500 -521
rect 1505 -525 1509 -521
rect 1515 -525 1519 -521
rect 1523 -525 1527 -521
rect 1532 -525 1536 -521
rect 1541 -525 1545 -521
rect 1550 -525 1554 -521
rect 1566 -525 1570 -521
rect 1575 -525 1579 -521
rect 1726 -531 1730 -527
rect 1950 -531 1954 -527
rect 1726 -540 1730 -536
rect 1950 -540 1954 -536
rect 1726 -549 1730 -545
rect 1950 -549 1954 -545
rect 1726 -558 1730 -554
rect 1950 -558 1954 -554
rect 1726 -566 1730 -562
rect 1950 -566 1954 -562
rect 1726 -576 1730 -572
rect 1950 -576 1954 -572
rect 1726 -585 1730 -581
rect 1950 -585 1954 -581
rect 1726 -594 1730 -590
rect 1950 -594 1954 -590
rect 1726 -602 1730 -598
rect 1950 -602 1954 -598
rect 1726 -612 1730 -608
rect 1950 -612 1954 -608
rect 1726 -621 1730 -617
rect 1950 -621 1954 -617
rect 1726 -648 1730 -644
rect 1950 -648 1954 -644
rect 1726 -657 1730 -653
rect 1950 -657 1954 -653
rect 1726 -666 1730 -662
rect 2972 -660 2976 -656
rect 2980 -660 2984 -656
rect 2989 -660 2993 -656
rect 2998 -660 3002 -656
rect 3008 -660 3012 -656
rect 3016 -660 3020 -656
rect 3025 -660 3029 -656
rect 3034 -660 3038 -656
rect 3061 -660 3065 -656
rect 3070 -660 3074 -656
rect 3080 -660 3084 -656
rect 3088 -660 3092 -656
rect 3097 -660 3101 -656
rect 3106 -660 3110 -656
rect 3116 -660 3120 -656
rect 3124 -660 3128 -656
rect 1950 -666 1954 -662
rect 3133 -660 3137 -656
rect 3142 -660 3146 -656
rect 3169 -660 3173 -656
rect 3178 -660 3182 -656
rect 3188 -660 3192 -656
rect 3196 -660 3200 -656
rect 1726 -674 1730 -670
rect 1950 -674 1954 -670
rect 3205 -660 3209 -656
rect 3214 -660 3218 -656
rect 3241 -660 3245 -656
rect 3250 -660 3254 -656
rect 3260 -660 3264 -656
rect 3268 -660 3272 -656
rect 3277 -660 3281 -656
rect 3286 -660 3290 -656
rect 3296 -660 3300 -656
rect 3304 -660 3308 -656
rect 3320 -660 3324 -656
rect 3329 -660 3333 -656
rect 1726 -684 1730 -680
rect 1950 -684 1954 -680
rect 1726 -693 1730 -689
rect 1950 -693 1954 -689
rect 1726 -720 1730 -716
rect 1950 -720 1954 -716
rect 1726 -729 1730 -725
rect 1950 -729 1954 -725
rect 1726 -738 1730 -734
rect 1950 -738 1954 -734
rect 1726 -746 1730 -742
rect 1950 -746 1954 -742
rect 1726 -756 1730 -752
rect 1950 -756 1954 -752
rect 1726 -765 1730 -761
rect 1726 -774 1730 -770
rect 1950 -765 1954 -761
rect 1950 -774 1954 -770
rect 1726 -782 1730 -778
rect 1950 -782 1954 -778
rect 1726 -792 1730 -788
rect 1950 -792 1954 -788
rect 1726 -801 1730 -797
rect 1950 -801 1954 -797
rect 1726 -828 1730 -824
rect 1950 -828 1954 -824
rect 1726 -837 1730 -833
rect 1950 -837 1954 -833
rect 1726 -846 1730 -842
rect 1950 -846 1954 -842
rect 1726 -854 1730 -850
rect 1950 -854 1954 -850
rect 1726 -864 1730 -860
rect 1950 -864 1954 -860
rect 1726 -873 1730 -869
rect 1950 -873 1954 -869
rect 1726 -882 1730 -878
rect 1950 -882 1954 -878
rect 1726 -890 1730 -886
rect 1950 -890 1954 -886
<< polysilicon >>
rect 1753 500 1756 502
rect 1776 501 1812 502
rect 1776 500 1819 501
rect 1912 501 1948 502
rect 1905 500 1948 501
rect 1968 500 1971 502
rect 1753 464 1756 466
rect 1776 465 1812 466
rect 1776 464 1819 465
rect 1912 465 1948 466
rect 1905 464 1948 465
rect 1968 464 1971 466
rect 1753 427 1789 429
rect 1799 427 1815 429
rect 1909 427 1925 429
rect 1935 427 1971 429
rect 1753 392 1756 394
rect 1776 392 1815 394
rect 1909 392 1948 394
rect 1968 392 1971 394
rect 1742 357 1789 358
rect 1736 356 1789 357
rect 1799 356 1817 358
rect 1907 356 1925 358
rect 1935 357 1982 358
rect 1935 356 1988 357
rect 1753 320 1789 322
rect 1799 320 1813 322
rect 3131 325 3132 331
rect 1911 320 1925 322
rect 1935 320 1971 322
rect 2986 311 2988 314
rect 3022 311 3024 314
rect 1741 284 1756 286
rect 1776 284 1817 286
rect 1907 284 1948 286
rect 1968 284 1983 286
rect 2986 255 2988 291
rect 3022 255 3024 291
rect 3059 278 3061 314
rect 3094 311 3096 314
rect 1754 248 1789 250
rect 1799 248 1813 250
rect 1911 248 1925 250
rect 1935 248 1970 250
rect 2987 248 2988 255
rect 3023 248 3024 255
rect 3059 252 3061 268
rect 3094 252 3096 291
rect 3130 278 3132 325
rect 3166 278 3168 314
rect 3202 311 3204 326
rect 3130 250 3132 268
rect 3166 254 3168 268
rect 3202 250 3204 291
rect 3238 278 3240 313
rect 3274 278 3276 325
rect 3310 311 3312 325
rect 3326 311 3328 322
rect 3310 278 3312 291
rect 3326 278 3328 291
rect 3238 254 3240 268
rect 3274 249 3276 268
rect 3310 248 3312 268
rect 3326 258 3328 268
rect 1742 212 1789 214
rect 1799 212 1818 214
rect 1906 212 1925 214
rect 1935 212 1982 214
rect 1742 176 1756 178
rect 1776 176 1789 178
rect 1799 176 1819 178
rect 1905 176 1925 178
rect 1935 176 1948 178
rect 1968 176 1982 178
rect 1745 158 1756 160
rect 1776 158 1789 160
rect 1799 158 1814 160
rect 1910 158 1925 160
rect 1935 158 1948 160
rect 1968 158 1979 160
rect 2987 150 2988 157
rect 3023 150 3024 157
rect 1745 142 1756 144
rect 1776 142 1789 144
rect 1799 142 1814 144
rect 1910 142 1925 144
rect 1935 142 1948 144
rect 1968 142 1979 144
rect 1355 130 1356 136
rect 1210 116 1212 119
rect 1246 116 1248 119
rect 1210 60 1212 96
rect 1246 60 1248 96
rect 1283 83 1285 119
rect 1318 116 1320 119
rect 1211 53 1212 60
rect 1247 53 1248 60
rect 1283 57 1285 73
rect 1318 57 1320 96
rect 1354 83 1356 130
rect 1390 83 1392 119
rect 1426 116 1428 131
rect 1354 55 1356 73
rect 1390 59 1392 73
rect 1426 55 1428 96
rect 1462 83 1464 118
rect 1498 83 1500 130
rect 1534 116 1536 130
rect 1552 116 1554 127
rect 1568 116 1570 127
rect 2986 114 2988 150
rect 3022 114 3024 150
rect 3059 137 3061 153
rect 1534 83 1536 96
rect 1552 83 1554 96
rect 1568 83 1570 96
rect 2986 91 2988 94
rect 3022 91 3024 94
rect 3059 91 3061 127
rect 3094 114 3096 153
rect 3130 137 3132 155
rect 3166 137 3168 151
rect 3094 91 3096 94
rect 3130 80 3132 127
rect 3166 91 3168 127
rect 3202 114 3204 155
rect 3238 137 3240 151
rect 3274 137 3276 156
rect 3310 137 3312 157
rect 3329 137 3331 147
rect 3131 74 3132 80
rect 3202 79 3204 94
rect 3238 92 3240 127
rect 3274 80 3276 127
rect 3310 114 3312 127
rect 3329 114 3331 127
rect 3310 80 3312 94
rect 3329 83 3331 94
rect 1462 59 1464 73
rect 1498 54 1500 73
rect 1534 53 1536 73
rect 1552 58 1554 73
rect 1568 58 1570 73
rect 2541 3 2543 6
rect 2557 3 2559 6
rect 2455 -7 2467 -6
rect 2455 -8 2457 -7
rect 2462 -8 2467 -7
rect 2517 -8 2521 -6
rect 1211 -27 1212 -20
rect 1247 -27 1248 -20
rect 1210 -63 1212 -27
rect 1246 -63 1248 -27
rect 1283 -40 1285 -24
rect 1210 -86 1212 -83
rect 1246 -86 1248 -83
rect 1283 -86 1285 -50
rect 1318 -63 1320 -24
rect 1354 -40 1356 -22
rect 1390 -40 1392 -26
rect 1318 -86 1320 -83
rect 1354 -97 1356 -50
rect 1390 -86 1392 -50
rect 1426 -63 1428 -22
rect 1462 -40 1464 -26
rect 1498 -40 1500 -21
rect 1534 -40 1536 -20
rect 2463 -24 2467 -22
rect 2517 -24 2521 -22
rect 1552 -40 1554 -25
rect 1568 -40 1570 -25
rect 2463 -30 2465 -24
rect 2541 -25 2543 -17
rect 2557 -25 2559 -17
rect 2542 -29 2543 -25
rect 2558 -29 2559 -25
rect 1712 -34 1714 -32
rect 1800 -34 1802 -32
rect 1889 -34 1891 -32
rect 1977 -34 1979 -32
rect 1712 -39 1713 -34
rect 1712 -44 1714 -39
rect 1728 -41 1736 -40
rect 1800 -39 1801 -34
rect 1741 -41 1747 -40
rect 1728 -42 1747 -41
rect 1757 -42 1761 -40
rect 1728 -44 1730 -42
rect 1355 -103 1356 -97
rect 1426 -98 1428 -83
rect 1462 -85 1464 -50
rect 1498 -97 1500 -50
rect 1534 -63 1536 -50
rect 1552 -63 1554 -50
rect 1568 -63 1570 -50
rect 1534 -97 1536 -83
rect 1552 -94 1554 -83
rect 1568 -94 1570 -83
rect 1800 -44 1802 -39
rect 1816 -41 1824 -40
rect 1889 -39 1890 -34
rect 1829 -41 1835 -40
rect 1816 -42 1835 -41
rect 1845 -42 1849 -40
rect 1816 -44 1818 -42
rect 1889 -44 1891 -39
rect 1905 -41 1913 -40
rect 1977 -39 1978 -34
rect 1918 -41 1924 -40
rect 1905 -42 1924 -41
rect 1934 -42 1938 -40
rect 1905 -44 1907 -42
rect 1977 -44 1979 -39
rect 1993 -41 2001 -40
rect 2464 -35 2465 -30
rect 2541 -32 2543 -29
rect 2557 -32 2559 -29
rect 2172 -38 2208 -36
rect 2228 -38 2262 -36
rect 2282 -38 2287 -36
rect 2006 -41 2012 -40
rect 1993 -42 2012 -41
rect 2022 -42 2026 -40
rect 1993 -44 1995 -42
rect 2463 -41 2465 -35
rect 2178 -50 2208 -48
rect 2228 -50 2262 -48
rect 2282 -50 2287 -48
rect 2541 -46 2543 -42
rect 2557 -46 2559 -42
rect 2463 -55 2465 -51
rect 2197 -68 2208 -66
rect 2228 -68 2252 -66
rect 2282 -68 2285 -66
rect 2204 -80 2208 -78
rect 2228 -80 2252 -78
rect 2282 -80 2284 -78
rect 2204 -92 2208 -90
rect 2228 -92 2252 -90
rect 2282 -92 2285 -90
rect 1712 -98 1714 -94
rect 1728 -98 1730 -94
rect 1800 -98 1802 -94
rect 1816 -98 1818 -94
rect 1889 -98 1891 -94
rect 1905 -98 1907 -94
rect 1977 -98 1979 -94
rect 1993 -98 1995 -94
rect 2037 -99 2042 -97
rect 2062 -99 2097 -97
rect 2117 -99 2120 -97
rect 2037 -111 2042 -109
rect 2062 -111 2097 -109
rect 2117 -111 2120 -109
rect 1700 -120 1703 -118
rect 1723 -119 1731 -118
rect 1735 -119 1738 -118
rect 1723 -120 1738 -119
rect 1748 -120 1752 -118
rect 1788 -120 1791 -118
rect 1811 -119 1819 -118
rect 1823 -119 1826 -118
rect 1811 -120 1826 -119
rect 1836 -120 1840 -118
rect 1877 -120 1880 -118
rect 1900 -119 1908 -118
rect 1912 -119 1915 -118
rect 1900 -120 1915 -119
rect 1925 -120 1929 -118
rect 1965 -120 1968 -118
rect 1988 -119 1996 -118
rect 2205 -116 2208 -114
rect 2228 -116 2252 -114
rect 2282 -116 2285 -114
rect 2290 -116 2293 -114
rect 2323 -116 2346 -114
rect 2366 -116 2369 -114
rect 2000 -119 2003 -118
rect 1988 -120 2003 -119
rect 2013 -120 2017 -118
rect 2037 -128 2042 -126
rect 2062 -128 2097 -126
rect 2117 -128 2120 -126
rect 2135 -128 2140 -126
rect 2160 -128 2178 -126
rect 2198 -128 2201 -126
rect 2205 -128 2208 -126
rect 2228 -128 2252 -126
rect 2282 -128 2285 -126
rect 2290 -128 2293 -126
rect 2323 -128 2346 -126
rect 2366 -128 2369 -126
rect 1700 -136 1703 -134
rect 1723 -135 1731 -134
rect 1735 -135 1738 -134
rect 1723 -136 1738 -135
rect 1748 -136 1752 -134
rect 1788 -136 1791 -134
rect 1811 -135 1819 -134
rect 1823 -135 1826 -134
rect 1811 -136 1826 -135
rect 1836 -136 1840 -134
rect 1877 -136 1880 -134
rect 1900 -135 1908 -134
rect 1912 -135 1915 -134
rect 1900 -136 1915 -135
rect 1925 -136 1929 -134
rect 1965 -136 1968 -134
rect 1988 -135 1996 -134
rect 2000 -135 2003 -134
rect 1988 -136 2003 -135
rect 2013 -136 2017 -134
rect 2986 -131 2987 -124
rect 3022 -131 3023 -124
rect 2037 -140 2042 -138
rect 2062 -140 2097 -138
rect 2117 -140 2120 -138
rect 2134 -140 2140 -138
rect 2160 -140 2178 -138
rect 2198 -140 2208 -138
rect 2228 -140 2252 -138
rect 2282 -140 2293 -138
rect 2323 -140 2346 -138
rect 2366 -140 2403 -138
rect 2985 -167 2987 -131
rect 3021 -167 3023 -131
rect 3058 -144 3060 -128
rect 2541 -183 2543 -180
rect 2557 -183 2559 -180
rect 2455 -193 2467 -192
rect 2455 -194 2457 -193
rect 2462 -194 2467 -193
rect 2517 -194 2521 -192
rect 2985 -190 2987 -187
rect 3021 -190 3023 -187
rect 3058 -190 3060 -154
rect 3093 -167 3095 -128
rect 3129 -144 3131 -126
rect 3165 -144 3167 -130
rect 3093 -190 3095 -187
rect 3129 -201 3131 -154
rect 3165 -190 3167 -154
rect 3201 -167 3203 -126
rect 3237 -144 3239 -130
rect 3273 -144 3275 -125
rect 3309 -144 3311 -124
rect 3326 -144 3328 -134
rect 2463 -210 2467 -208
rect 2517 -210 2521 -208
rect 2463 -216 2465 -210
rect 2541 -211 2543 -203
rect 2557 -211 2559 -203
rect 3130 -207 3131 -201
rect 3201 -202 3203 -187
rect 3237 -189 3239 -154
rect 3273 -201 3275 -154
rect 3309 -167 3311 -154
rect 3326 -167 3328 -154
rect 3309 -201 3311 -187
rect 3326 -198 3328 -187
rect 2542 -215 2543 -211
rect 2558 -215 2559 -211
rect 2464 -221 2465 -216
rect 2541 -218 2543 -215
rect 2557 -218 2559 -215
rect 2463 -227 2465 -221
rect 2541 -232 2543 -228
rect 2557 -232 2559 -228
rect 2463 -241 2465 -237
rect 1350 -291 1351 -285
rect 1205 -305 1207 -302
rect 1241 -305 1243 -302
rect 1205 -361 1207 -325
rect 1241 -361 1243 -325
rect 1278 -338 1280 -302
rect 1313 -305 1315 -302
rect 1206 -368 1207 -361
rect 1242 -368 1243 -361
rect 1278 -364 1280 -348
rect 1313 -364 1315 -325
rect 1349 -338 1351 -291
rect 1385 -338 1387 -302
rect 1421 -305 1423 -290
rect 1703 -290 1705 -285
rect 1715 -290 1717 -285
rect 1759 -290 1761 -285
rect 1771 -290 1773 -285
rect 1812 -290 1814 -285
rect 1824 -290 1826 -285
rect 1868 -290 1870 -285
rect 1880 -290 1882 -285
rect 1349 -366 1351 -348
rect 1385 -362 1387 -348
rect 1421 -366 1423 -325
rect 1457 -338 1459 -303
rect 1493 -338 1495 -291
rect 1529 -305 1531 -291
rect 1547 -305 1549 -294
rect 1563 -305 1565 -294
rect 1529 -338 1531 -325
rect 1547 -338 1549 -325
rect 1563 -338 1565 -325
rect 1703 -336 1705 -310
rect 1715 -336 1717 -310
rect 1739 -311 1741 -308
rect 1739 -336 1741 -321
rect 1759 -336 1761 -310
rect 1771 -336 1773 -310
rect 1795 -311 1797 -308
rect 1795 -336 1797 -321
rect 1812 -336 1814 -310
rect 1824 -336 1826 -310
rect 1847 -311 1849 -308
rect 1847 -336 1849 -321
rect 1868 -336 1870 -310
rect 1880 -336 1882 -310
rect 1903 -311 1905 -308
rect 1923 -311 1925 -308
rect 1941 -311 1943 -308
rect 1970 -316 1973 -314
rect 1993 -316 2031 -314
rect 2071 -316 2078 -314
rect 1903 -336 1905 -321
rect 1923 -336 1925 -321
rect 1941 -336 1943 -321
rect 1958 -328 1973 -326
rect 1993 -328 2031 -326
rect 2071 -328 2074 -326
rect 1457 -362 1459 -348
rect 1493 -367 1495 -348
rect 1529 -368 1531 -348
rect 1547 -363 1549 -348
rect 1563 -363 1565 -348
rect 1970 -340 1973 -338
rect 1993 -339 2015 -338
rect 2020 -339 2031 -338
rect 1993 -340 2031 -339
rect 2071 -340 2074 -338
rect 1970 -352 1973 -350
rect 1993 -352 2031 -350
rect 2071 -352 2074 -350
rect 1703 -366 1705 -356
rect 1704 -368 1705 -366
rect 1715 -367 1717 -356
rect 1739 -359 1741 -356
rect 1759 -366 1761 -356
rect 1771 -366 1773 -356
rect 1795 -359 1797 -356
rect 1812 -366 1814 -356
rect 1824 -366 1826 -356
rect 1847 -359 1849 -356
rect 1868 -366 1870 -356
rect 1880 -366 1882 -356
rect 1903 -359 1905 -356
rect 1923 -359 1925 -356
rect 1941 -359 1943 -356
rect 1970 -370 1973 -368
rect 1993 -370 2031 -368
rect 2071 -370 2078 -368
rect 1970 -382 1973 -380
rect 1993 -382 2031 -380
rect 2071 -382 2074 -380
rect 1970 -394 1973 -392
rect 1993 -394 2031 -392
rect 2071 -394 2073 -392
rect 2541 -398 2543 -395
rect 2557 -398 2559 -395
rect 1970 -406 1973 -404
rect 1993 -406 2031 -404
rect 2071 -406 2073 -404
rect 2455 -408 2467 -407
rect 2455 -409 2457 -408
rect 2462 -409 2467 -408
rect 2517 -409 2521 -407
rect 2463 -425 2467 -423
rect 2517 -425 2521 -423
rect 2463 -431 2465 -425
rect 2541 -426 2543 -418
rect 2557 -426 2559 -418
rect 3131 -421 3132 -415
rect 2542 -430 2543 -426
rect 2558 -430 2559 -426
rect 2464 -436 2465 -431
rect 2541 -433 2543 -430
rect 2557 -433 2559 -430
rect 2463 -442 2465 -436
rect 1206 -461 1207 -454
rect 1242 -461 1243 -454
rect 2986 -435 2988 -432
rect 3022 -435 3024 -432
rect 2541 -447 2543 -443
rect 2557 -447 2559 -443
rect 1205 -497 1207 -461
rect 1241 -497 1243 -461
rect 1278 -474 1280 -458
rect 1205 -520 1207 -517
rect 1241 -520 1243 -517
rect 1278 -520 1280 -484
rect 1313 -497 1315 -458
rect 1349 -474 1351 -456
rect 1385 -474 1387 -460
rect 1313 -520 1315 -517
rect 1349 -531 1351 -484
rect 1385 -520 1387 -484
rect 1421 -497 1423 -456
rect 1457 -474 1459 -460
rect 1493 -474 1495 -455
rect 1529 -474 1531 -454
rect 2463 -456 2465 -452
rect 1547 -474 1549 -459
rect 1563 -474 1565 -459
rect 1350 -537 1351 -531
rect 1421 -532 1423 -517
rect 1457 -519 1459 -484
rect 1493 -531 1495 -484
rect 1529 -497 1531 -484
rect 1547 -497 1549 -484
rect 1563 -497 1565 -484
rect 2986 -491 2988 -455
rect 3022 -491 3024 -455
rect 3059 -468 3061 -432
rect 3094 -435 3096 -432
rect 2987 -498 2988 -491
rect 3023 -498 3024 -491
rect 3059 -494 3061 -478
rect 3094 -494 3096 -455
rect 3130 -468 3132 -421
rect 3166 -468 3168 -432
rect 3202 -435 3204 -420
rect 3130 -496 3132 -478
rect 3166 -492 3168 -478
rect 3202 -496 3204 -455
rect 3238 -468 3240 -433
rect 3274 -468 3276 -421
rect 3310 -435 3312 -421
rect 3326 -435 3328 -424
rect 3310 -468 3312 -455
rect 3326 -468 3328 -455
rect 3238 -492 3240 -478
rect 3274 -497 3276 -478
rect 3310 -498 3312 -478
rect 3326 -488 3328 -478
rect 1529 -531 1531 -517
rect 1547 -528 1549 -517
rect 1563 -528 1565 -517
rect 1723 -518 1734 -516
rect 1754 -518 1767 -516
rect 1777 -518 1792 -516
rect 1888 -518 1903 -516
rect 1913 -518 1926 -516
rect 1946 -518 1957 -516
rect 1723 -534 1734 -532
rect 1754 -534 1767 -532
rect 1777 -534 1792 -532
rect 1888 -534 1903 -532
rect 1913 -534 1926 -532
rect 1946 -534 1957 -532
rect 1720 -552 1734 -550
rect 1754 -552 1767 -550
rect 1777 -552 1797 -550
rect 1883 -552 1903 -550
rect 1913 -552 1926 -550
rect 1946 -552 1960 -550
rect 1720 -588 1767 -586
rect 1777 -588 1796 -586
rect 1884 -588 1903 -586
rect 1913 -588 1960 -586
rect 2987 -596 2988 -589
rect 3023 -596 3024 -589
rect 1732 -624 1767 -622
rect 1777 -624 1791 -622
rect 1889 -624 1903 -622
rect 1913 -624 1948 -622
rect 2986 -632 2988 -596
rect 3022 -632 3024 -596
rect 3059 -609 3061 -593
rect 2986 -655 2988 -652
rect 3022 -655 3024 -652
rect 3059 -655 3061 -619
rect 3094 -632 3096 -593
rect 3130 -609 3132 -591
rect 3166 -609 3168 -595
rect 3094 -655 3096 -652
rect 1719 -660 1734 -658
rect 1754 -660 1795 -658
rect 1885 -660 1926 -658
rect 1946 -660 1961 -658
rect 3130 -666 3132 -619
rect 3166 -655 3168 -619
rect 3202 -632 3204 -591
rect 3238 -609 3240 -595
rect 3274 -609 3276 -590
rect 3310 -609 3312 -589
rect 3326 -609 3328 -599
rect 3131 -672 3132 -666
rect 3202 -667 3204 -652
rect 3238 -654 3240 -619
rect 3274 -666 3276 -619
rect 3310 -632 3312 -619
rect 3326 -632 3328 -619
rect 3310 -666 3312 -652
rect 3326 -663 3328 -652
rect 1731 -696 1767 -694
rect 1777 -696 1791 -694
rect 1889 -696 1903 -694
rect 1913 -696 1949 -694
rect 1714 -731 1767 -730
rect 1720 -732 1767 -731
rect 1777 -732 1795 -730
rect 1885 -732 1903 -730
rect 1913 -731 1966 -730
rect 1913 -732 1960 -731
rect 1731 -768 1734 -766
rect 1754 -768 1793 -766
rect 1887 -768 1926 -766
rect 1946 -768 1949 -766
rect 1731 -803 1767 -801
rect 1777 -803 1793 -801
rect 1887 -803 1903 -801
rect 1913 -803 1949 -801
rect 1731 -840 1734 -838
rect 1754 -839 1797 -838
rect 1754 -840 1790 -839
rect 1883 -839 1926 -838
rect 1890 -840 1926 -839
rect 1946 -840 1949 -838
rect 1731 -876 1734 -874
rect 1754 -875 1797 -874
rect 1754 -876 1790 -875
rect 1883 -875 1926 -874
rect 1890 -876 1926 -875
rect 1946 -876 1949 -874
<< polycontact >>
rect 1812 501 1819 508
rect 1905 501 1912 508
rect 1815 424 1822 431
rect 1902 424 1909 431
rect 1736 357 1742 363
rect 1982 357 1988 363
rect 3125 325 3131 331
rect 3200 326 3206 333
rect 1734 282 1741 288
rect 1983 282 1990 288
rect 2980 248 2987 255
rect 3272 325 3278 331
rect 3305 325 3315 333
rect 3057 245 3064 252
rect 3321 281 3326 286
rect 1736 210 1742 216
rect 1982 210 1988 216
rect 1734 173 1742 183
rect 1982 173 1990 183
rect 1780 160 1785 165
rect 1939 160 1944 165
rect 2980 150 2987 157
rect 3057 153 3064 160
rect 1780 144 1785 148
rect 1939 144 1944 148
rect 1349 130 1355 136
rect 1424 131 1430 138
rect 1204 53 1211 60
rect 1496 130 1502 136
rect 1529 130 1539 138
rect 1281 50 1288 57
rect 1547 87 1552 92
rect 1564 87 1568 92
rect 3125 74 3131 80
rect 3324 119 3329 124
rect 3200 72 3206 79
rect 3272 74 3278 80
rect 3305 72 3315 80
rect 2457 -12 2462 -7
rect 1204 -27 1211 -20
rect 1281 -24 1288 -17
rect 2538 -29 2542 -25
rect 2554 -29 2558 -25
rect 1713 -39 1718 -34
rect 1736 -41 1741 -36
rect 1801 -39 1806 -34
rect 1349 -103 1355 -97
rect 1547 -59 1552 -54
rect 1564 -59 1568 -54
rect 1824 -41 1829 -36
rect 1890 -39 1895 -34
rect 1913 -41 1918 -36
rect 1978 -39 1983 -34
rect 2001 -41 2006 -36
rect 2459 -35 2464 -30
rect 2192 -71 2197 -66
rect 1424 -105 1430 -98
rect 1496 -103 1502 -97
rect 1529 -105 1539 -97
rect 2236 -97 2241 -92
rect 1731 -119 1735 -115
rect 1819 -119 1823 -115
rect 1908 -119 1912 -115
rect 1996 -119 2000 -115
rect 2085 -116 2090 -111
rect 1731 -135 1735 -131
rect 1819 -135 1823 -131
rect 1908 -135 1912 -131
rect 1996 -135 2000 -131
rect 2979 -131 2986 -124
rect 3056 -128 3063 -121
rect 2403 -142 2408 -137
rect 2457 -198 2462 -193
rect 3124 -207 3130 -201
rect 3321 -162 3326 -157
rect 3199 -209 3205 -202
rect 3271 -207 3277 -201
rect 3304 -209 3314 -201
rect 2538 -215 2542 -211
rect 2554 -215 2558 -211
rect 2459 -221 2464 -216
rect 1344 -291 1350 -285
rect 1419 -290 1425 -283
rect 1199 -368 1206 -361
rect 1491 -291 1497 -285
rect 1524 -291 1534 -283
rect 1276 -371 1283 -364
rect 1542 -334 1547 -329
rect 1559 -334 1563 -329
rect 1734 -332 1739 -327
rect 1790 -332 1795 -327
rect 1842 -332 1847 -327
rect 1898 -332 1903 -327
rect 1919 -328 1923 -324
rect 1937 -328 1941 -324
rect 1953 -329 1958 -324
rect 2016 -380 2021 -375
rect 2073 -396 2078 -391
rect 2073 -407 2077 -403
rect 2457 -413 2462 -408
rect 3125 -421 3131 -415
rect 3200 -420 3206 -413
rect 2538 -430 2542 -426
rect 2554 -430 2558 -426
rect 2459 -436 2464 -431
rect 1199 -461 1206 -454
rect 1276 -458 1283 -451
rect 1344 -537 1350 -531
rect 1542 -493 1547 -488
rect 1559 -493 1563 -488
rect 2980 -498 2987 -491
rect 3272 -421 3278 -415
rect 3305 -421 3315 -413
rect 3057 -501 3064 -494
rect 3321 -465 3326 -460
rect 1758 -522 1763 -518
rect 1917 -522 1922 -518
rect 1419 -539 1425 -532
rect 1491 -537 1497 -531
rect 1524 -539 1534 -531
rect 1758 -539 1763 -534
rect 1917 -539 1922 -534
rect 1712 -557 1720 -547
rect 1960 -557 1968 -547
rect 1714 -590 1720 -584
rect 1960 -590 1966 -584
rect 2980 -596 2987 -589
rect 3057 -593 3064 -586
rect 1712 -662 1719 -656
rect 1961 -662 1968 -656
rect 3125 -672 3131 -666
rect 3321 -627 3326 -622
rect 3200 -674 3206 -667
rect 3272 -672 3278 -666
rect 3305 -674 3315 -666
rect 1714 -737 1720 -731
rect 1960 -737 1966 -731
rect 1793 -805 1800 -798
rect 1880 -805 1887 -798
rect 1790 -882 1797 -875
rect 1883 -882 1890 -875
<< metal1 >>
rect 1745 549 1979 552
rect 1745 519 1748 549
rect 1976 519 1979 549
rect 1745 516 1752 519
rect 1745 512 1748 516
rect 1745 508 1752 512
rect 1745 504 1748 508
rect 1801 517 1809 519
rect 1801 513 1803 517
rect 1807 513 1809 517
rect 1801 508 1809 513
rect 1752 504 1756 507
rect 1745 503 1756 504
rect 1801 504 1803 508
rect 1807 504 1809 508
rect 1745 499 1752 503
rect 1745 495 1748 499
rect 1745 490 1752 495
rect 1745 486 1748 490
rect 1745 480 1752 486
rect 1745 476 1748 480
rect 1745 472 1752 476
rect 1745 468 1748 472
rect 1745 463 1752 468
rect 1756 471 1776 495
rect 1801 491 1809 504
rect 1812 512 1830 519
rect 1812 508 1819 512
rect 1801 487 1803 491
rect 1807 487 1809 491
rect 1801 481 1809 487
rect 1801 477 1803 481
rect 1807 477 1809 481
rect 1801 472 1809 477
rect 1801 468 1803 472
rect 1807 468 1809 472
rect 1745 459 1748 463
rect 1745 454 1752 459
rect 1745 450 1748 454
rect 1727 288 1733 367
rect 1736 363 1742 430
rect 1745 427 1752 450
rect 1756 439 1776 459
rect 1762 434 1776 439
rect 1801 455 1809 468
rect 1801 451 1803 455
rect 1807 451 1809 455
rect 1801 445 1809 451
rect 1801 441 1803 445
rect 1807 441 1809 445
rect 1801 436 1809 441
rect 1762 430 1789 434
rect 1801 432 1803 436
rect 1807 432 1809 436
rect 1745 423 1748 427
rect 1801 426 1809 432
rect 1823 431 1830 512
rect 1745 418 1752 423
rect 1799 422 1809 426
rect 1822 424 1830 431
rect 1894 512 1912 519
rect 1894 431 1901 512
rect 1905 508 1912 512
rect 1915 517 1923 519
rect 1915 513 1917 517
rect 1921 513 1923 517
rect 1915 508 1923 513
rect 1915 504 1917 508
rect 1921 504 1923 508
rect 1972 516 1979 519
rect 1976 512 1979 516
rect 1972 508 1979 512
rect 1915 491 1923 504
rect 1968 504 1972 507
rect 1976 504 1979 508
rect 1968 503 1979 504
rect 1972 499 1979 503
rect 1915 487 1917 491
rect 1921 487 1923 491
rect 1915 481 1923 487
rect 1915 477 1917 481
rect 1921 477 1923 481
rect 1915 472 1923 477
rect 1915 468 1917 472
rect 1921 468 1923 472
rect 1915 455 1923 468
rect 1948 471 1968 495
rect 1976 495 1979 499
rect 1972 490 1979 495
rect 1976 486 1979 490
rect 1972 480 1979 486
rect 1976 476 1979 480
rect 1972 472 1979 476
rect 1976 468 1979 472
rect 1972 463 1979 468
rect 1915 451 1917 455
rect 1921 451 1923 455
rect 1915 445 1923 451
rect 1915 441 1917 445
rect 1921 441 1923 445
rect 1915 436 1923 441
rect 1915 432 1917 436
rect 1921 432 1923 436
rect 1948 439 1968 459
rect 1948 434 1962 439
rect 1894 424 1902 431
rect 1915 426 1923 432
rect 1935 430 1962 434
rect 1976 459 1979 463
rect 1972 454 1979 459
rect 1976 450 1979 454
rect 1972 427 1979 450
rect 1745 414 1748 418
rect 1745 408 1752 414
rect 1745 404 1748 408
rect 1745 400 1752 404
rect 1745 396 1748 400
rect 1801 419 1809 422
rect 1801 415 1803 419
rect 1807 415 1809 419
rect 1801 409 1809 415
rect 1801 405 1803 409
rect 1807 405 1809 409
rect 1801 400 1809 405
rect 1752 396 1756 399
rect 1745 395 1756 396
rect 1801 396 1803 400
rect 1807 396 1809 400
rect 1915 422 1925 426
rect 1976 423 1979 427
rect 1915 419 1923 422
rect 1915 415 1917 419
rect 1921 415 1923 419
rect 1915 409 1923 415
rect 1915 405 1917 409
rect 1921 405 1923 409
rect 1915 400 1923 405
rect 1915 396 1917 400
rect 1921 396 1923 400
rect 1972 418 1979 423
rect 1976 414 1979 418
rect 1972 408 1979 414
rect 1976 404 1979 408
rect 1972 400 1979 404
rect 1745 391 1752 395
rect 1745 387 1748 391
rect 1745 382 1752 387
rect 1745 378 1748 382
rect 1745 372 1752 378
rect 1745 368 1748 372
rect 1745 364 1752 368
rect 1745 360 1748 364
rect 1745 355 1752 360
rect 1756 375 1776 387
rect 1762 367 1776 375
rect 1756 363 1776 367
rect 1801 383 1809 396
rect 1801 379 1803 383
rect 1807 380 1809 383
rect 1915 383 1923 396
rect 1968 396 1972 399
rect 1976 396 1979 400
rect 1968 395 1979 396
rect 1972 391 1979 395
rect 1915 380 1917 383
rect 1807 379 1858 380
rect 1801 377 1858 379
rect 1801 373 1809 377
rect 1863 379 1917 380
rect 1921 379 1923 383
rect 1863 377 1923 379
rect 1801 369 1803 373
rect 1807 369 1809 373
rect 1801 364 1809 369
rect 1756 359 1789 363
rect 1801 360 1803 364
rect 1807 360 1809 364
rect 1745 351 1748 355
rect 1745 346 1752 351
rect 1745 342 1748 346
rect 1745 319 1752 342
rect 1789 327 1798 351
rect 1801 347 1809 360
rect 1801 343 1803 347
rect 1807 343 1809 347
rect 1801 337 1809 343
rect 1801 333 1803 337
rect 1807 333 1809 337
rect 1801 328 1809 333
rect 1801 324 1803 328
rect 1807 324 1809 328
rect 1915 373 1923 377
rect 1915 369 1917 373
rect 1921 369 1923 373
rect 1915 364 1923 369
rect 1915 360 1917 364
rect 1921 360 1923 364
rect 1948 375 1968 387
rect 1948 367 1962 375
rect 1948 363 1968 367
rect 1915 347 1923 360
rect 1935 359 1968 363
rect 1976 387 1979 391
rect 1972 382 1979 387
rect 1976 378 1979 382
rect 1972 372 1979 378
rect 1976 368 1979 372
rect 1972 364 1979 368
rect 1976 360 1979 364
rect 1972 355 1979 360
rect 1982 363 1988 430
rect 1915 343 1917 347
rect 1921 343 1923 347
rect 1915 337 1923 343
rect 1915 333 1917 337
rect 1921 333 1923 337
rect 1915 328 1923 333
rect 1915 324 1917 328
rect 1921 324 1923 328
rect 1801 319 1809 324
rect 1745 315 1748 319
rect 1799 315 1809 319
rect 1915 319 1923 324
rect 1926 327 1935 351
rect 1976 351 1979 355
rect 1972 346 1979 351
rect 1976 342 1979 346
rect 1972 319 1979 342
rect 1745 310 1752 315
rect 1745 306 1748 310
rect 1745 300 1752 306
rect 1745 296 1748 300
rect 1745 292 1752 296
rect 1745 288 1748 292
rect 1801 311 1809 315
rect 1801 307 1803 311
rect 1807 307 1809 311
rect 1801 301 1809 307
rect 1801 297 1803 301
rect 1807 297 1809 301
rect 1801 292 1809 297
rect 1752 288 1756 291
rect 1727 282 1734 288
rect 1745 287 1756 288
rect 1801 288 1803 292
rect 1807 288 1809 292
rect 1745 283 1752 287
rect 1727 216 1733 282
rect 1745 279 1748 283
rect 1745 274 1752 279
rect 1745 270 1748 274
rect 1745 247 1752 270
rect 1756 261 1776 279
rect 1763 255 1776 261
rect 1801 275 1809 288
rect 1801 271 1803 275
rect 1807 271 1809 275
rect 1801 265 1809 271
rect 1801 261 1803 265
rect 1807 261 1809 265
rect 1801 256 1809 261
rect 1763 251 1789 255
rect 1801 252 1803 256
rect 1807 252 1809 256
rect 1915 315 1925 319
rect 1976 315 1979 319
rect 1915 311 1923 315
rect 1915 307 1917 311
rect 1921 307 1923 311
rect 1915 301 1923 307
rect 1915 297 1917 301
rect 1921 297 1923 301
rect 1915 292 1923 297
rect 1915 288 1917 292
rect 1921 288 1923 292
rect 1972 310 1979 315
rect 1976 306 1979 310
rect 1972 300 1979 306
rect 1976 296 1979 300
rect 1972 292 1979 296
rect 1915 275 1923 288
rect 1968 288 1972 291
rect 1976 288 1979 292
rect 1991 288 1997 367
rect 3121 334 3278 340
rect 3200 333 3206 334
rect 3058 325 3125 331
rect 3272 331 3278 334
rect 3305 333 3315 342
rect 2969 319 3373 322
rect 2969 315 2972 319
rect 2976 315 2980 319
rect 2984 315 2989 319
rect 2993 315 2998 319
rect 3002 315 3008 319
rect 3012 315 3016 319
rect 3020 315 3025 319
rect 3029 315 3034 319
rect 3038 315 3061 319
rect 3065 315 3070 319
rect 3074 315 3080 319
rect 3084 315 3088 319
rect 3092 315 3097 319
rect 3101 315 3106 319
rect 3110 315 3116 319
rect 3120 315 3124 319
rect 3128 315 3133 319
rect 3137 315 3142 319
rect 3146 315 3169 319
rect 3173 315 3178 319
rect 3182 315 3188 319
rect 3192 315 3196 319
rect 3200 315 3205 319
rect 3209 315 3214 319
rect 3218 315 3241 319
rect 3245 315 3250 319
rect 3254 315 3260 319
rect 3264 315 3268 319
rect 3272 315 3277 319
rect 3281 315 3286 319
rect 3290 315 3296 319
rect 3300 315 3304 319
rect 3308 315 3329 319
rect 3333 318 3373 319
rect 3333 315 3339 318
rect 2981 311 2985 315
rect 3089 311 3093 315
rect 3197 311 3201 315
rect 3305 311 3309 315
rect 3321 311 3325 315
rect 2993 291 3017 311
rect 3029 305 3049 311
rect 3029 291 3058 305
rect 3101 305 3113 311
rect 3121 305 3129 311
rect 3101 291 3129 305
rect 3209 304 3227 311
rect 3209 291 3237 304
rect 1968 287 1979 288
rect 1972 283 1979 287
rect 1915 271 1917 275
rect 1921 271 1923 275
rect 1915 265 1923 271
rect 1915 261 1917 265
rect 1921 261 1923 265
rect 1915 256 1923 261
rect 1915 252 1917 256
rect 1921 252 1923 256
rect 1948 261 1968 279
rect 1948 255 1961 261
rect 1745 243 1748 247
rect 1745 238 1752 243
rect 1745 234 1748 238
rect 1745 228 1752 234
rect 1745 224 1748 228
rect 1745 220 1752 224
rect 1745 216 1748 220
rect 1727 210 1736 216
rect 1745 211 1752 216
rect 1789 219 1798 243
rect 1801 239 1809 252
rect 1801 235 1803 239
rect 1807 235 1809 239
rect 1801 229 1809 235
rect 1801 225 1803 229
rect 1807 225 1809 229
rect 1801 220 1809 225
rect 1801 216 1803 220
rect 1807 216 1809 220
rect 1801 211 1809 216
rect 1745 207 1748 211
rect 1799 207 1809 211
rect 1745 202 1752 207
rect 1745 198 1748 202
rect 1745 192 1752 198
rect 1745 188 1748 192
rect 1745 184 1752 188
rect 1725 173 1734 183
rect 1745 180 1748 184
rect 1801 203 1809 207
rect 1801 199 1803 203
rect 1807 199 1809 203
rect 1801 193 1809 199
rect 1801 189 1803 193
rect 1807 189 1809 193
rect 1801 184 1809 189
rect 1801 183 1803 184
rect 1752 180 1756 183
rect 1745 179 1756 180
rect 1799 180 1803 183
rect 1807 180 1809 184
rect 1799 179 1809 180
rect 1745 175 1752 179
rect 1745 171 1748 175
rect 1776 171 1789 175
rect 1745 166 1752 171
rect 1745 162 1748 166
rect 1780 165 1785 171
rect 1801 166 1809 179
rect 1801 165 1803 166
rect 1752 162 1756 165
rect 1745 161 1756 162
rect 1745 157 1752 161
rect 1799 162 1803 165
rect 1807 162 1809 166
rect 1799 161 1809 162
rect 1345 139 1502 145
rect 1424 138 1430 139
rect 1282 130 1349 136
rect 1496 136 1502 139
rect 1529 138 1539 147
rect 1745 153 1748 157
rect 1776 153 1789 157
rect 1745 149 1752 153
rect 1745 145 1756 149
rect 1780 148 1785 153
rect 1801 150 1809 161
rect 1801 149 1803 150
rect 1745 141 1752 145
rect 1799 146 1803 149
rect 1807 146 1809 150
rect 1799 145 1809 146
rect 1745 137 1748 141
rect 1776 137 1789 141
rect 1745 132 1752 137
rect 1745 128 1748 132
rect 1745 127 1752 128
rect 1160 125 1752 127
rect 1160 124 1748 125
rect 1160 122 1196 124
rect 1160 -91 1163 122
rect 1193 120 1196 122
rect 1200 120 1204 124
rect 1208 120 1213 124
rect 1217 120 1222 124
rect 1226 120 1232 124
rect 1236 120 1240 124
rect 1244 120 1249 124
rect 1253 120 1258 124
rect 1262 120 1285 124
rect 1289 120 1294 124
rect 1298 120 1304 124
rect 1308 120 1312 124
rect 1316 120 1321 124
rect 1325 120 1330 124
rect 1334 120 1340 124
rect 1344 120 1348 124
rect 1352 120 1357 124
rect 1361 120 1366 124
rect 1370 120 1393 124
rect 1397 120 1402 124
rect 1406 120 1412 124
rect 1416 120 1420 124
rect 1424 120 1429 124
rect 1433 120 1438 124
rect 1442 120 1465 124
rect 1469 120 1474 124
rect 1478 120 1484 124
rect 1488 120 1492 124
rect 1496 120 1501 124
rect 1505 120 1510 124
rect 1514 120 1520 124
rect 1524 120 1528 124
rect 1532 120 1537 124
rect 1541 120 1546 124
rect 1550 120 1555 124
rect 1559 120 1571 124
rect 1575 120 1580 124
rect 1584 123 1748 124
rect 1584 120 1587 123
rect 1205 116 1209 120
rect 1313 116 1317 120
rect 1421 116 1425 120
rect 1529 116 1533 120
rect 1547 116 1551 120
rect 1563 116 1567 120
rect 1217 96 1241 116
rect 1253 110 1273 116
rect 1253 96 1282 110
rect 1325 110 1337 116
rect 1345 110 1353 116
rect 1325 96 1353 110
rect 1433 109 1451 116
rect 1433 96 1461 109
rect 1278 83 1282 96
rect 1349 83 1353 96
rect 1457 83 1461 96
rect 1537 92 1541 96
rect 1555 92 1559 96
rect 1537 87 1547 92
rect 1555 87 1564 92
rect 1571 90 1575 96
rect 1537 83 1541 87
rect 1555 83 1559 87
rect 1571 85 1766 90
rect 1571 83 1575 85
rect 1361 74 1385 83
rect 1286 71 1290 73
rect 1469 74 1493 83
rect 1393 71 1397 73
rect 1501 71 1505 73
rect 1529 71 1533 73
rect 1547 71 1551 73
rect 1563 71 1567 73
rect 1193 69 1587 71
rect 1193 65 1195 69
rect 1199 65 1204 69
rect 1208 65 1221 69
rect 1225 65 1231 69
rect 1235 65 1240 69
rect 1244 65 1257 69
rect 1261 65 1267 69
rect 1271 65 1276 69
rect 1280 65 1293 69
rect 1297 65 1303 69
rect 1307 65 1312 69
rect 1316 65 1329 69
rect 1333 65 1339 69
rect 1343 65 1348 69
rect 1352 65 1365 69
rect 1369 65 1375 69
rect 1379 65 1384 69
rect 1388 65 1401 69
rect 1405 65 1411 69
rect 1415 65 1420 69
rect 1424 65 1437 69
rect 1441 65 1447 69
rect 1451 65 1456 69
rect 1460 65 1473 69
rect 1477 65 1483 69
rect 1487 65 1492 69
rect 1496 65 1509 69
rect 1513 65 1519 69
rect 1523 65 1528 69
rect 1532 65 1546 69
rect 1550 65 1562 69
rect 1566 65 1579 69
rect 1583 65 1587 69
rect 1193 63 1587 65
rect 1193 53 1204 60
rect 1193 49 1200 53
rect 1281 49 1288 50
rect 1193 42 1288 49
rect 1330 20 1333 63
rect 1193 -16 1288 -9
rect 1193 -20 1200 -16
rect 1281 -17 1288 -16
rect 1193 -27 1204 -20
rect 1330 -30 1333 15
rect 1761 9 1766 85
rect 1781 36 1786 137
rect 1801 133 1809 145
rect 1801 129 1803 133
rect 1807 129 1809 133
rect 1801 125 1809 129
rect 1915 239 1923 252
rect 1935 251 1961 255
rect 1976 279 1979 283
rect 1990 282 1997 288
rect 1972 274 1979 279
rect 1976 270 1979 274
rect 1972 247 1979 270
rect 1915 235 1917 239
rect 1921 235 1923 239
rect 1915 229 1923 235
rect 1915 225 1917 229
rect 1921 225 1923 229
rect 1915 220 1923 225
rect 1915 216 1917 220
rect 1921 216 1923 220
rect 1915 211 1923 216
rect 1926 219 1935 243
rect 1976 243 1979 247
rect 1972 238 1979 243
rect 1976 234 1979 238
rect 1972 228 1979 234
rect 1976 224 1979 228
rect 1972 220 1979 224
rect 1976 216 1979 220
rect 1991 216 1997 282
rect 3054 278 3058 291
rect 3125 278 3129 291
rect 3233 278 3237 291
rect 3313 286 3317 291
rect 3313 281 3321 286
rect 3329 284 3333 291
rect 3313 278 3317 281
rect 3329 279 3336 284
rect 3329 278 3333 279
rect 3137 269 3161 278
rect 3062 266 3066 268
rect 3245 269 3269 278
rect 3169 266 3173 268
rect 3277 266 3281 268
rect 3305 266 3309 268
rect 3321 266 3325 268
rect 2969 264 3339 266
rect 2969 260 2971 264
rect 2975 260 2980 264
rect 2984 260 2997 264
rect 3001 260 3007 264
rect 3011 260 3016 264
rect 3020 260 3033 264
rect 3037 260 3043 264
rect 3047 260 3052 264
rect 3056 260 3069 264
rect 3073 260 3079 264
rect 3083 260 3088 264
rect 3092 260 3105 264
rect 3109 260 3115 264
rect 3119 260 3124 264
rect 3128 260 3141 264
rect 3145 260 3151 264
rect 3155 260 3160 264
rect 3164 260 3177 264
rect 3181 260 3187 264
rect 3191 260 3196 264
rect 3200 260 3213 264
rect 3217 260 3223 264
rect 3227 260 3232 264
rect 3236 260 3249 264
rect 3253 260 3259 264
rect 3263 260 3268 264
rect 3272 260 3285 264
rect 3289 260 3295 264
rect 3299 260 3304 264
rect 3308 260 3320 264
rect 3324 260 3339 264
rect 2969 258 3339 260
rect 2969 248 2980 255
rect 2969 244 2976 248
rect 3057 244 3064 245
rect 2969 242 3064 244
rect 1972 211 1979 216
rect 1915 207 1925 211
rect 1976 207 1979 211
rect 1988 210 1997 216
rect 2708 237 3064 242
rect 1915 203 1923 207
rect 1915 199 1917 203
rect 1921 199 1923 203
rect 1915 193 1923 199
rect 1915 189 1917 193
rect 1921 189 1923 193
rect 1915 184 1923 189
rect 1915 180 1917 184
rect 1921 183 1923 184
rect 1972 202 1979 207
rect 1976 198 1979 202
rect 1972 192 1979 198
rect 1976 188 1979 192
rect 1972 184 1979 188
rect 1921 180 1925 183
rect 1915 179 1925 180
rect 1968 180 1972 183
rect 1976 180 1979 184
rect 1968 179 1979 180
rect 1915 166 1923 179
rect 1972 175 1979 179
rect 1935 171 1948 175
rect 1976 171 1979 175
rect 1990 173 1999 183
rect 1915 162 1917 166
rect 1921 165 1923 166
rect 1939 165 1944 171
rect 1972 166 1979 171
rect 1921 162 1925 165
rect 1915 161 1925 162
rect 1915 150 1923 161
rect 1968 162 1972 165
rect 1976 162 1979 166
rect 1968 161 1979 162
rect 1972 157 1979 161
rect 1935 153 1948 157
rect 1976 153 1979 157
rect 1915 146 1917 150
rect 1921 149 1923 150
rect 1921 146 1925 149
rect 1915 145 1925 146
rect 1939 148 1944 153
rect 1972 149 1979 153
rect 1915 133 1923 145
rect 1968 145 1979 149
rect 1972 141 1979 145
rect 1935 137 1948 141
rect 1976 137 1979 141
rect 1915 129 1917 133
rect 1921 129 1923 133
rect 1915 125 1923 129
rect 1939 45 1944 137
rect 1972 132 1979 137
rect 1976 128 1979 132
rect 1972 125 1979 128
rect 1975 -10 1979 125
rect 2182 12 2570 15
rect 2182 -10 2185 12
rect 2433 10 2532 12
rect 2433 9 2437 10
rect 1691 -14 2390 -10
rect 1193 -32 1587 -30
rect 1193 -36 1195 -32
rect 1199 -36 1204 -32
rect 1208 -36 1221 -32
rect 1225 -36 1231 -32
rect 1235 -36 1240 -32
rect 1244 -36 1257 -32
rect 1261 -36 1267 -32
rect 1271 -36 1276 -32
rect 1280 -36 1293 -32
rect 1297 -36 1303 -32
rect 1307 -36 1312 -32
rect 1316 -36 1329 -32
rect 1333 -36 1339 -32
rect 1343 -36 1348 -32
rect 1352 -36 1365 -32
rect 1369 -36 1375 -32
rect 1379 -36 1384 -32
rect 1388 -36 1401 -32
rect 1405 -36 1411 -32
rect 1415 -36 1420 -32
rect 1424 -36 1437 -32
rect 1441 -36 1447 -32
rect 1451 -36 1456 -32
rect 1460 -36 1473 -32
rect 1477 -36 1483 -32
rect 1487 -36 1492 -32
rect 1496 -36 1509 -32
rect 1513 -36 1519 -32
rect 1523 -36 1528 -32
rect 1532 -36 1546 -32
rect 1550 -36 1562 -32
rect 1566 -36 1579 -32
rect 1583 -36 1587 -32
rect 1193 -38 1587 -36
rect 1286 -40 1290 -38
rect 1393 -40 1397 -38
rect 1361 -50 1385 -41
rect 1501 -40 1505 -38
rect 1469 -50 1493 -41
rect 1529 -40 1533 -38
rect 1547 -40 1551 -38
rect 1563 -40 1567 -38
rect 1278 -63 1282 -50
rect 1349 -63 1353 -50
rect 1457 -63 1461 -50
rect 1537 -54 1541 -50
rect 1555 -54 1559 -50
rect 1537 -59 1547 -54
rect 1555 -59 1564 -54
rect 1571 -55 1659 -50
rect 1537 -63 1541 -59
rect 1555 -63 1559 -59
rect 1571 -63 1575 -55
rect 1217 -83 1241 -63
rect 1253 -77 1282 -63
rect 1253 -83 1273 -77
rect 1325 -77 1353 -63
rect 1325 -83 1337 -77
rect 1345 -83 1353 -77
rect 1433 -76 1461 -63
rect 1433 -83 1451 -76
rect 1205 -87 1209 -83
rect 1313 -87 1317 -83
rect 1421 -87 1425 -83
rect 1529 -87 1533 -83
rect 1547 -87 1551 -83
rect 1563 -87 1567 -83
rect 1193 -91 1196 -87
rect 1200 -91 1204 -87
rect 1208 -91 1213 -87
rect 1217 -91 1222 -87
rect 1226 -91 1232 -87
rect 1236 -91 1240 -87
rect 1244 -91 1249 -87
rect 1253 -91 1258 -87
rect 1262 -91 1285 -87
rect 1289 -91 1294 -87
rect 1298 -91 1304 -87
rect 1308 -91 1312 -87
rect 1316 -91 1321 -87
rect 1325 -91 1330 -87
rect 1334 -91 1340 -87
rect 1344 -91 1348 -87
rect 1352 -91 1357 -87
rect 1361 -91 1366 -87
rect 1370 -91 1393 -87
rect 1397 -91 1402 -87
rect 1406 -91 1412 -87
rect 1416 -91 1420 -87
rect 1424 -91 1429 -87
rect 1433 -91 1438 -87
rect 1442 -91 1465 -87
rect 1469 -91 1474 -87
rect 1478 -91 1484 -87
rect 1488 -91 1492 -87
rect 1496 -91 1501 -87
rect 1505 -91 1510 -87
rect 1514 -91 1520 -87
rect 1524 -91 1528 -87
rect 1532 -91 1537 -87
rect 1541 -91 1546 -87
rect 1550 -91 1555 -87
rect 1559 -91 1571 -87
rect 1575 -91 1580 -87
rect 1584 -91 1587 -87
rect 1160 -94 1587 -91
rect 1169 -294 1172 -94
rect 1282 -103 1349 -97
rect 1424 -106 1430 -105
rect 1496 -106 1502 -103
rect 1345 -112 1502 -106
rect 1529 -114 1539 -105
rect 1691 -106 1694 -14
rect 1747 -25 1770 -18
rect 1707 -30 1731 -25
rect 1707 -31 1711 -30
rect 1707 -42 1710 -31
rect 1718 -39 1722 -34
rect 1707 -44 1711 -42
rect 1723 -44 1727 -39
rect 1736 -36 1741 -25
rect 1747 -35 1757 -25
rect 1715 -102 1719 -94
rect 1731 -102 1735 -94
rect 1747 -102 1757 -47
rect 1715 -106 1757 -102
rect 1691 -109 1699 -106
rect 1691 -113 1694 -109
rect 1698 -113 1699 -109
rect 1691 -117 1703 -113
rect 1731 -115 1735 -106
rect 1764 -113 1770 -25
rect 1691 -124 1699 -117
rect 1748 -117 1770 -113
rect 1691 -128 1694 -124
rect 1698 -128 1699 -124
rect 1723 -122 1728 -121
rect 1723 -125 1740 -122
rect 1691 -129 1699 -128
rect 1691 -133 1703 -129
rect 1731 -131 1735 -125
rect 1764 -129 1770 -117
rect 1691 -139 1699 -133
rect 1748 -133 1770 -129
rect 1691 -143 1694 -139
rect 1698 -143 1699 -139
rect 1723 -138 1728 -137
rect 1723 -141 1740 -138
rect 1691 -147 1699 -143
rect 1691 -148 1696 -147
rect 1340 -282 1497 -276
rect 1419 -283 1425 -282
rect 1277 -291 1344 -285
rect 1491 -285 1497 -282
rect 1524 -283 1534 -274
rect 1169 -297 1582 -294
rect 1169 -299 1191 -297
rect 1169 -523 1174 -299
rect 1188 -301 1191 -299
rect 1195 -301 1199 -297
rect 1203 -301 1208 -297
rect 1212 -301 1217 -297
rect 1221 -301 1227 -297
rect 1231 -301 1235 -297
rect 1239 -301 1244 -297
rect 1248 -301 1253 -297
rect 1257 -301 1280 -297
rect 1284 -301 1289 -297
rect 1293 -301 1299 -297
rect 1303 -301 1307 -297
rect 1311 -301 1316 -297
rect 1320 -301 1325 -297
rect 1329 -301 1335 -297
rect 1339 -301 1343 -297
rect 1347 -301 1352 -297
rect 1356 -301 1361 -297
rect 1365 -301 1388 -297
rect 1392 -301 1397 -297
rect 1401 -301 1407 -297
rect 1411 -301 1415 -297
rect 1419 -301 1424 -297
rect 1428 -301 1433 -297
rect 1437 -301 1460 -297
rect 1464 -301 1469 -297
rect 1473 -301 1479 -297
rect 1483 -301 1487 -297
rect 1491 -301 1496 -297
rect 1500 -301 1505 -297
rect 1509 -301 1515 -297
rect 1519 -301 1523 -297
rect 1527 -301 1532 -297
rect 1536 -301 1541 -297
rect 1545 -301 1550 -297
rect 1554 -301 1566 -297
rect 1570 -301 1575 -297
rect 1579 -301 1582 -297
rect 1200 -305 1204 -301
rect 1308 -305 1312 -301
rect 1416 -305 1420 -301
rect 1524 -305 1528 -301
rect 1542 -305 1546 -301
rect 1558 -305 1562 -301
rect 1212 -325 1236 -305
rect 1248 -311 1268 -305
rect 1248 -325 1277 -311
rect 1320 -311 1332 -305
rect 1340 -311 1348 -305
rect 1320 -325 1348 -311
rect 1428 -312 1446 -305
rect 1428 -325 1456 -312
rect 1273 -338 1277 -325
rect 1344 -338 1348 -325
rect 1452 -338 1456 -325
rect 1532 -329 1536 -325
rect 1550 -329 1554 -325
rect 1532 -334 1542 -329
rect 1550 -334 1559 -329
rect 1566 -331 1570 -325
rect 1532 -338 1536 -334
rect 1550 -338 1554 -334
rect 1566 -336 1677 -331
rect 1566 -338 1570 -336
rect 1356 -347 1380 -338
rect 1281 -350 1285 -348
rect 1464 -347 1488 -338
rect 1388 -350 1392 -348
rect 1496 -350 1500 -348
rect 1524 -350 1528 -348
rect 1542 -350 1546 -348
rect 1558 -350 1562 -348
rect 1188 -352 1582 -350
rect 1188 -356 1190 -352
rect 1194 -356 1199 -352
rect 1203 -356 1216 -352
rect 1220 -356 1226 -352
rect 1230 -356 1235 -352
rect 1239 -356 1252 -352
rect 1256 -356 1262 -352
rect 1266 -356 1271 -352
rect 1275 -356 1288 -352
rect 1292 -356 1298 -352
rect 1302 -356 1307 -352
rect 1311 -356 1324 -352
rect 1328 -356 1334 -352
rect 1338 -356 1343 -352
rect 1347 -356 1360 -352
rect 1364 -356 1370 -352
rect 1374 -356 1379 -352
rect 1383 -356 1396 -352
rect 1400 -356 1406 -352
rect 1410 -356 1415 -352
rect 1419 -356 1432 -352
rect 1436 -356 1442 -352
rect 1446 -356 1451 -352
rect 1455 -356 1468 -352
rect 1472 -356 1478 -352
rect 1482 -356 1487 -352
rect 1491 -356 1504 -352
rect 1508 -356 1514 -352
rect 1518 -356 1523 -352
rect 1527 -356 1541 -352
rect 1545 -356 1557 -352
rect 1561 -356 1574 -352
rect 1578 -356 1582 -352
rect 1188 -358 1582 -356
rect 1188 -368 1199 -361
rect 1188 -372 1195 -368
rect 1276 -372 1283 -371
rect 1188 -379 1283 -372
rect 1394 -408 1399 -358
rect 1691 -360 1694 -148
rect 1731 -205 1736 -141
rect 1764 -151 1770 -133
rect 1779 -106 1784 -14
rect 1835 -25 1858 -18
rect 1795 -30 1819 -25
rect 1795 -31 1799 -30
rect 1795 -42 1798 -31
rect 1806 -39 1810 -34
rect 1795 -44 1799 -42
rect 1811 -44 1815 -39
rect 1824 -36 1829 -25
rect 1835 -35 1845 -25
rect 1803 -102 1807 -94
rect 1819 -102 1823 -94
rect 1835 -102 1845 -47
rect 1803 -106 1845 -102
rect 1779 -109 1787 -106
rect 1779 -113 1782 -109
rect 1786 -113 1787 -109
rect 1779 -117 1791 -113
rect 1819 -115 1823 -106
rect 1852 -113 1858 -25
rect 1779 -122 1787 -117
rect 1836 -117 1858 -113
rect 1779 -126 1782 -122
rect 1786 -126 1787 -122
rect 1811 -122 1816 -121
rect 1811 -125 1828 -122
rect 1779 -129 1787 -126
rect 1779 -133 1791 -129
rect 1819 -131 1823 -125
rect 1852 -129 1858 -117
rect 1779 -138 1787 -133
rect 1836 -133 1858 -129
rect 1779 -142 1782 -138
rect 1786 -142 1787 -138
rect 1811 -138 1816 -137
rect 1811 -141 1828 -138
rect 1779 -147 1787 -142
rect 1819 -197 1824 -141
rect 1852 -151 1858 -133
rect 1868 -106 1873 -14
rect 1924 -25 1947 -18
rect 1884 -30 1908 -25
rect 1884 -31 1888 -30
rect 1884 -42 1887 -31
rect 1895 -39 1899 -34
rect 1884 -44 1888 -42
rect 1900 -44 1904 -39
rect 1913 -36 1918 -25
rect 1924 -35 1934 -25
rect 1892 -102 1896 -94
rect 1908 -102 1912 -94
rect 1924 -102 1934 -47
rect 1892 -106 1934 -102
rect 1868 -109 1876 -106
rect 1868 -113 1871 -109
rect 1875 -113 1876 -109
rect 1868 -117 1880 -113
rect 1908 -115 1912 -106
rect 1941 -113 1947 -25
rect 1868 -129 1876 -117
rect 1925 -117 1947 -113
rect 1900 -122 1905 -121
rect 1900 -125 1917 -122
rect 1868 -133 1871 -129
rect 1875 -133 1880 -129
rect 1908 -131 1912 -125
rect 1941 -129 1947 -117
rect 1868 -140 1876 -133
rect 1925 -133 1947 -129
rect 1868 -144 1871 -140
rect 1875 -144 1876 -140
rect 1900 -138 1905 -137
rect 1900 -141 1917 -138
rect 1868 -147 1876 -144
rect 1908 -189 1912 -141
rect 1941 -151 1947 -133
rect 1956 -106 1961 -14
rect 2012 -25 2035 -18
rect 1972 -30 1996 -25
rect 1972 -31 1976 -30
rect 1972 -42 1975 -31
rect 1983 -39 1987 -34
rect 1972 -44 1976 -42
rect 1988 -44 1992 -39
rect 2001 -36 2006 -25
rect 2012 -35 2022 -25
rect 1980 -102 1984 -94
rect 1996 -102 2000 -94
rect 2012 -102 2022 -47
rect 1980 -106 2022 -102
rect 1956 -109 1964 -106
rect 1956 -113 1959 -109
rect 1963 -113 1964 -109
rect 1956 -117 1968 -113
rect 1996 -115 2000 -106
rect 2029 -112 2035 -25
rect 2062 -96 2073 -92
rect 2120 -92 2124 -14
rect 2202 -15 2390 -14
rect 2078 -96 2093 -92
rect 2117 -96 2124 -92
rect 2088 -102 2093 -96
rect 2088 -106 2097 -102
rect 2029 -113 2042 -112
rect 1956 -124 1964 -117
rect 2013 -116 2042 -113
rect 2120 -112 2124 -96
rect 2117 -116 2124 -112
rect 2013 -117 2035 -116
rect 1956 -128 1959 -124
rect 1963 -128 1964 -124
rect 1988 -122 1993 -121
rect 1988 -125 2005 -122
rect 1956 -129 1964 -128
rect 1956 -133 1968 -129
rect 1996 -131 2000 -125
rect 2029 -129 2035 -117
rect 2085 -121 2090 -116
rect 2120 -121 2124 -116
rect 2062 -125 2093 -121
rect 2117 -125 2124 -121
rect 1956 -140 1964 -133
rect 2013 -133 2035 -129
rect 2088 -131 2093 -125
rect 1956 -144 1959 -140
rect 1963 -144 1964 -140
rect 1988 -138 1993 -137
rect 1988 -141 2005 -138
rect 2029 -141 2035 -133
rect 2088 -135 2097 -131
rect 1956 -147 1964 -144
rect 1956 -157 1961 -147
rect 1996 -163 2001 -141
rect 2029 -145 2042 -141
rect 2120 -141 2124 -125
rect 2117 -145 2124 -141
rect 2129 -141 2134 -26
rect 2202 -31 2205 -15
rect 2202 -35 2208 -31
rect 2231 -35 2262 -31
rect 2202 -51 2205 -35
rect 2231 -41 2236 -35
rect 2228 -45 2236 -41
rect 2202 -55 2208 -51
rect 2163 -71 2192 -66
rect 2202 -71 2205 -55
rect 2228 -65 2242 -61
rect 2247 -65 2252 -61
rect 2163 -121 2168 -71
rect 2202 -75 2208 -71
rect 2202 -93 2205 -75
rect 2228 -87 2232 -65
rect 2202 -97 2208 -93
rect 2202 -119 2205 -97
rect 2236 -109 2241 -97
rect 2262 -98 2267 -35
rect 2282 -55 2296 -51
rect 2292 -93 2296 -55
rect 2282 -97 2296 -93
rect 2228 -113 2252 -109
rect 2202 -121 2208 -119
rect 2160 -125 2174 -121
rect 2198 -123 2208 -121
rect 2198 -125 2205 -123
rect 2169 -131 2174 -125
rect 2169 -135 2178 -131
rect 2202 -141 2205 -125
rect 2228 -135 2232 -113
rect 2287 -141 2290 -97
rect 2323 -113 2346 -109
rect 2129 -145 2140 -141
rect 2198 -145 2208 -141
rect 2282 -145 2293 -141
rect 2029 -151 2035 -145
rect 2129 -151 2134 -145
rect 2202 -146 2205 -145
rect 2287 -151 2290 -145
rect 2035 -156 2290 -151
rect 2342 -152 2346 -113
rect 2385 -119 2390 -15
rect 2366 -123 2390 -119
rect 2385 -141 2390 -123
rect 2366 -145 2390 -141
rect 2403 -137 2408 -30
rect 2342 -155 2344 -152
rect 1996 -168 2381 -163
rect 1908 -194 2006 -189
rect 2011 -194 2085 -189
rect 2090 -194 2235 -189
rect 2240 -193 2365 -189
rect 2403 -197 2408 -142
rect 1819 -202 2015 -197
rect 2020 -202 2408 -197
rect 2433 -171 2436 9
rect 2529 8 2532 10
rect 2536 8 2545 12
rect 2549 8 2561 12
rect 2565 8 2570 12
rect 2529 7 2570 8
rect 2536 3 2540 7
rect 2552 3 2556 7
rect 2448 -4 2467 -1
rect 2448 -5 2454 -4
rect 2465 -5 2467 -4
rect 2448 -25 2453 -5
rect 2457 -16 2462 -12
rect 2517 -13 2529 -9
rect 2462 -21 2467 -17
rect 2525 -25 2529 -13
rect 2544 -22 2548 -17
rect 2560 -22 2564 -17
rect 2545 -25 2548 -22
rect 2561 -25 2564 -22
rect 2708 -25 2713 237
rect 3184 209 3188 258
rect 2517 -29 2538 -25
rect 2545 -29 2554 -25
rect 2448 -35 2459 -30
rect 2525 -41 2529 -29
rect 2441 -51 2458 -41
rect 2470 -51 2529 -41
rect 2545 -34 2548 -29
rect 2561 -30 2713 -25
rect 2754 164 3064 168
rect 2561 -34 2564 -30
rect 2441 -58 2448 -51
rect 2536 -58 2540 -42
rect 2552 -58 2556 -42
rect 2441 -64 2574 -58
rect 2433 -174 2570 -171
rect 2433 -176 2532 -174
rect 2433 -177 2437 -176
rect 1731 -210 2025 -205
rect 2030 -210 2184 -205
rect 2189 -210 2334 -205
rect 2339 -210 2403 -205
rect 1725 -231 2085 -226
rect 2090 -231 2339 -226
rect 1718 -327 1722 -310
rect 1725 -327 1730 -231
rect 1742 -239 2047 -234
rect 1742 -315 1746 -239
rect 1781 -247 2290 -242
rect 1708 -332 1734 -327
rect 1708 -336 1712 -332
rect 1742 -336 1746 -321
rect 1774 -327 1778 -310
rect 1781 -327 1786 -247
rect 1798 -255 2172 -250
rect 1798 -315 1802 -255
rect 1827 -263 2064 -258
rect 1764 -332 1790 -327
rect 1764 -336 1768 -332
rect 1798 -336 1802 -321
rect 1827 -305 1832 -263
rect 1831 -306 1832 -305
rect 1850 -271 2161 -266
rect 2166 -271 2325 -266
rect 1827 -327 1831 -310
rect 1850 -315 1854 -271
rect 1883 -279 2046 -274
rect 1817 -332 1842 -327
rect 1817 -336 1821 -332
rect 1850 -336 1854 -321
rect 1883 -305 1887 -279
rect 1883 -327 1887 -310
rect 1944 -287 2075 -282
rect 2080 -287 2244 -282
rect 1906 -324 1910 -321
rect 1944 -315 1948 -287
rect 1964 -295 2071 -290
rect 2066 -301 2071 -295
rect 2412 -301 2416 -300
rect 2066 -305 2416 -301
rect 2066 -309 2071 -305
rect 1926 -324 1930 -321
rect 1944 -324 1948 -321
rect 1967 -313 1973 -309
rect 1873 -332 1898 -327
rect 1906 -328 1913 -324
rect 1873 -336 1877 -332
rect 1906 -336 1910 -328
rect 1918 -328 1919 -324
rect 1926 -328 1937 -324
rect 1926 -336 1930 -328
rect 1944 -329 1953 -324
rect 1944 -336 1948 -329
rect 1967 -331 1970 -313
rect 1993 -323 2002 -319
rect 1967 -335 1973 -331
rect 1698 -360 1702 -356
rect 1718 -360 1722 -356
rect 1734 -360 1738 -356
rect 1754 -360 1758 -356
rect 1774 -360 1778 -356
rect 1790 -360 1794 -356
rect 1807 -360 1811 -356
rect 1827 -360 1831 -356
rect 1842 -360 1846 -356
rect 1863 -360 1867 -356
rect 1883 -360 1887 -356
rect 1898 -360 1902 -356
rect 1918 -360 1922 -356
rect 1936 -360 1940 -356
rect 1967 -353 1970 -335
rect 1997 -343 2002 -323
rect 1993 -347 2002 -343
rect 1997 -353 2002 -347
rect 1967 -357 1973 -353
rect 1997 -357 2031 -353
rect 1967 -360 1970 -357
rect 1691 -363 1970 -360
rect 1967 -367 1973 -363
rect 1188 -450 1283 -443
rect 1188 -454 1195 -450
rect 1276 -451 1283 -450
rect 1188 -461 1199 -454
rect 1394 -464 1399 -413
rect 1188 -466 1582 -464
rect 1188 -470 1190 -466
rect 1194 -470 1199 -466
rect 1203 -470 1216 -466
rect 1220 -470 1226 -466
rect 1230 -470 1235 -466
rect 1239 -470 1252 -466
rect 1256 -470 1262 -466
rect 1266 -470 1271 -466
rect 1275 -470 1288 -466
rect 1292 -470 1298 -466
rect 1302 -470 1307 -466
rect 1311 -470 1324 -466
rect 1328 -470 1334 -466
rect 1338 -470 1343 -466
rect 1347 -470 1360 -466
rect 1364 -470 1370 -466
rect 1374 -470 1379 -466
rect 1383 -470 1396 -466
rect 1400 -470 1406 -466
rect 1410 -470 1415 -466
rect 1419 -470 1432 -466
rect 1436 -470 1442 -466
rect 1446 -470 1451 -466
rect 1455 -470 1468 -466
rect 1472 -470 1478 -466
rect 1482 -470 1487 -466
rect 1491 -470 1504 -466
rect 1508 -470 1514 -466
rect 1518 -470 1523 -466
rect 1527 -470 1541 -466
rect 1545 -470 1557 -466
rect 1561 -470 1574 -466
rect 1578 -470 1582 -466
rect 1188 -472 1582 -470
rect 1281 -474 1285 -472
rect 1388 -474 1392 -472
rect 1356 -484 1380 -475
rect 1496 -474 1500 -472
rect 1464 -484 1488 -475
rect 1524 -474 1528 -472
rect 1542 -474 1546 -472
rect 1558 -474 1562 -472
rect 1674 -484 1679 -380
rect 1967 -385 1970 -367
rect 1993 -377 2002 -373
rect 1967 -389 1973 -385
rect 1816 -397 1921 -392
rect 1273 -497 1277 -484
rect 1344 -497 1348 -484
rect 1452 -497 1456 -484
rect 1532 -488 1536 -484
rect 1550 -488 1554 -484
rect 1532 -493 1542 -488
rect 1550 -493 1559 -488
rect 1566 -489 1679 -484
rect 1532 -497 1536 -493
rect 1550 -497 1554 -493
rect 1566 -497 1570 -489
rect 1212 -517 1236 -497
rect 1248 -511 1277 -497
rect 1248 -517 1268 -511
rect 1320 -511 1348 -497
rect 1320 -517 1332 -511
rect 1340 -517 1348 -511
rect 1428 -510 1456 -497
rect 1428 -517 1446 -510
rect 1723 -502 1730 -499
rect 1723 -506 1726 -502
rect 1723 -511 1730 -506
rect 1758 -511 1763 -416
rect 1779 -503 1787 -499
rect 1779 -507 1781 -503
rect 1785 -507 1787 -503
rect 1723 -515 1726 -511
rect 1754 -515 1767 -511
rect 1200 -521 1204 -517
rect 1308 -521 1312 -517
rect 1416 -521 1420 -517
rect 1524 -521 1528 -517
rect 1542 -521 1546 -517
rect 1558 -521 1562 -517
rect 1723 -519 1730 -515
rect 1188 -523 1191 -521
rect 1169 -525 1191 -523
rect 1195 -525 1199 -521
rect 1203 -525 1208 -521
rect 1212 -525 1217 -521
rect 1221 -525 1227 -521
rect 1231 -525 1235 -521
rect 1239 -525 1244 -521
rect 1248 -525 1253 -521
rect 1257 -525 1280 -521
rect 1284 -525 1289 -521
rect 1293 -525 1299 -521
rect 1303 -525 1307 -521
rect 1311 -525 1316 -521
rect 1320 -525 1325 -521
rect 1329 -525 1335 -521
rect 1339 -525 1343 -521
rect 1347 -525 1352 -521
rect 1356 -525 1361 -521
rect 1365 -525 1388 -521
rect 1392 -525 1397 -521
rect 1401 -525 1407 -521
rect 1411 -525 1415 -521
rect 1419 -525 1424 -521
rect 1428 -525 1433 -521
rect 1437 -525 1460 -521
rect 1464 -525 1469 -521
rect 1473 -525 1479 -521
rect 1483 -525 1487 -521
rect 1491 -525 1496 -521
rect 1500 -525 1505 -521
rect 1509 -525 1515 -521
rect 1519 -525 1523 -521
rect 1527 -525 1532 -521
rect 1536 -525 1541 -521
rect 1545 -525 1550 -521
rect 1554 -525 1566 -521
rect 1570 -525 1575 -521
rect 1579 -525 1582 -521
rect 1169 -528 1582 -525
rect 1723 -523 1734 -519
rect 1779 -519 1787 -507
rect 1723 -527 1730 -523
rect 1758 -527 1763 -522
rect 1777 -520 1787 -519
rect 1777 -523 1781 -520
rect 1779 -524 1781 -523
rect 1785 -524 1787 -520
rect 1169 -905 1173 -528
rect 1723 -531 1726 -527
rect 1754 -531 1767 -527
rect 1277 -537 1344 -531
rect 1419 -540 1425 -539
rect 1491 -540 1497 -537
rect 1340 -546 1497 -540
rect 1524 -548 1534 -539
rect 1723 -535 1730 -531
rect 1723 -536 1734 -535
rect 1723 -540 1726 -536
rect 1730 -539 1734 -536
rect 1779 -535 1787 -524
rect 1777 -536 1787 -535
rect 1777 -539 1781 -536
rect 1723 -545 1730 -540
rect 1758 -545 1763 -539
rect 1779 -540 1781 -539
rect 1785 -540 1787 -536
rect 1703 -557 1712 -547
rect 1723 -549 1726 -545
rect 1754 -549 1767 -545
rect 1723 -553 1730 -549
rect 1779 -553 1787 -540
rect 1723 -554 1734 -553
rect 1723 -558 1726 -554
rect 1730 -557 1734 -554
rect 1777 -554 1787 -553
rect 1777 -557 1781 -554
rect 1723 -562 1730 -558
rect 1723 -566 1726 -562
rect 1723 -572 1730 -566
rect 1723 -576 1726 -572
rect 1723 -581 1730 -576
rect 1779 -558 1781 -557
rect 1785 -558 1787 -554
rect 1779 -563 1787 -558
rect 1779 -567 1781 -563
rect 1785 -567 1787 -563
rect 1779 -573 1787 -567
rect 1779 -577 1781 -573
rect 1785 -577 1787 -573
rect 1779 -581 1787 -577
rect 1705 -590 1714 -584
rect 1723 -585 1726 -581
rect 1777 -585 1787 -581
rect 1723 -590 1730 -585
rect 1705 -656 1711 -590
rect 1723 -594 1726 -590
rect 1723 -598 1730 -594
rect 1723 -602 1726 -598
rect 1723 -608 1730 -602
rect 1723 -612 1726 -608
rect 1723 -617 1730 -612
rect 1723 -621 1726 -617
rect 1767 -617 1776 -593
rect 1779 -590 1787 -585
rect 1779 -594 1781 -590
rect 1785 -594 1787 -590
rect 1779 -599 1787 -594
rect 1779 -603 1781 -599
rect 1785 -603 1787 -599
rect 1779 -609 1787 -603
rect 1779 -613 1781 -609
rect 1785 -613 1787 -609
rect 1723 -644 1730 -621
rect 1723 -648 1726 -644
rect 1723 -653 1730 -648
rect 1705 -662 1712 -656
rect 1723 -657 1726 -653
rect 1741 -629 1767 -625
rect 1779 -626 1787 -613
rect 1893 -503 1901 -499
rect 1893 -507 1895 -503
rect 1899 -507 1901 -503
rect 1893 -519 1901 -507
rect 1916 -511 1921 -397
rect 1967 -407 1970 -389
rect 1997 -397 2002 -377
rect 2016 -375 2021 -357
rect 2066 -363 2071 -313
rect 2078 -396 2262 -391
rect 1993 -401 2002 -397
rect 1997 -407 2002 -401
rect 2077 -407 2343 -403
rect 1967 -411 1973 -407
rect 1997 -411 2031 -407
rect 1950 -502 1957 -499
rect 1954 -506 1957 -502
rect 1950 -511 1957 -506
rect 1913 -515 1926 -511
rect 1954 -515 1957 -511
rect 1893 -520 1903 -519
rect 1893 -524 1895 -520
rect 1899 -523 1903 -520
rect 1950 -519 1957 -515
rect 1899 -524 1901 -523
rect 1893 -535 1901 -524
rect 1917 -527 1922 -522
rect 1946 -523 1957 -519
rect 1950 -527 1957 -523
rect 1913 -531 1926 -527
rect 1954 -531 1957 -527
rect 1893 -536 1903 -535
rect 1893 -540 1895 -536
rect 1899 -539 1903 -536
rect 1950 -535 1957 -531
rect 1946 -536 1957 -535
rect 1946 -539 1950 -536
rect 1899 -540 1901 -539
rect 1893 -553 1901 -540
rect 1917 -545 1922 -539
rect 1954 -540 1957 -536
rect 1950 -545 1957 -540
rect 1913 -549 1926 -545
rect 1954 -549 1957 -545
rect 1950 -553 1957 -549
rect 1893 -554 1903 -553
rect 1893 -558 1895 -554
rect 1899 -557 1903 -554
rect 1946 -554 1957 -553
rect 1946 -557 1950 -554
rect 1899 -558 1901 -557
rect 1893 -563 1901 -558
rect 1893 -567 1895 -563
rect 1899 -567 1901 -563
rect 1893 -573 1901 -567
rect 1893 -577 1895 -573
rect 1899 -577 1901 -573
rect 1893 -581 1901 -577
rect 1954 -558 1957 -554
rect 1968 -557 1977 -547
rect 1950 -562 1957 -558
rect 1954 -566 1957 -562
rect 1950 -572 1957 -566
rect 1954 -576 1957 -572
rect 1950 -581 1957 -576
rect 1893 -585 1903 -581
rect 1954 -585 1957 -581
rect 2013 -578 2018 -411
rect 2412 -462 2416 -305
rect 2433 -386 2436 -177
rect 2529 -178 2532 -176
rect 2536 -178 2545 -174
rect 2549 -178 2561 -174
rect 2565 -178 2570 -174
rect 2529 -179 2570 -178
rect 2536 -183 2540 -179
rect 2552 -183 2556 -179
rect 2448 -190 2467 -187
rect 2448 -191 2454 -190
rect 2465 -191 2467 -190
rect 2448 -211 2453 -191
rect 2457 -202 2462 -198
rect 2517 -199 2529 -195
rect 2462 -207 2467 -203
rect 2525 -211 2529 -199
rect 2544 -208 2548 -203
rect 2560 -208 2564 -203
rect 2545 -211 2548 -208
rect 2561 -211 2564 -208
rect 2754 -211 2759 164
rect 2969 161 3064 164
rect 2969 157 2976 161
rect 3057 160 3064 161
rect 2969 150 2980 157
rect 3184 147 3188 204
rect 2969 145 3348 147
rect 2969 141 2971 145
rect 2975 141 2980 145
rect 2984 141 2997 145
rect 3001 141 3007 145
rect 3011 141 3016 145
rect 3020 141 3033 145
rect 3037 141 3043 145
rect 3047 141 3052 145
rect 3056 141 3069 145
rect 3073 141 3079 145
rect 3083 141 3088 145
rect 3092 141 3105 145
rect 3109 141 3115 145
rect 3119 141 3124 145
rect 3128 141 3141 145
rect 3145 141 3151 145
rect 3155 141 3160 145
rect 3164 141 3177 145
rect 3181 141 3187 145
rect 3191 141 3196 145
rect 3200 141 3213 145
rect 3217 141 3223 145
rect 3227 141 3232 145
rect 3236 141 3249 145
rect 3253 141 3259 145
rect 3263 141 3268 145
rect 3272 141 3285 145
rect 3289 141 3295 145
rect 3299 141 3304 145
rect 3308 141 3323 145
rect 3327 141 3340 145
rect 3344 141 3348 145
rect 2969 139 3348 141
rect 3062 137 3066 139
rect 3169 137 3173 139
rect 3137 127 3161 136
rect 3277 137 3281 139
rect 3245 127 3269 136
rect 3305 137 3309 139
rect 3324 137 3328 139
rect 3054 114 3058 127
rect 3125 114 3129 127
rect 3233 114 3237 127
rect 3313 124 3317 127
rect 3332 126 3336 127
rect 3313 119 3324 124
rect 3332 121 3348 126
rect 3313 114 3317 119
rect 3332 114 3336 121
rect 2993 94 3017 114
rect 3029 100 3058 114
rect 3029 94 3049 100
rect 3101 100 3129 114
rect 3101 94 3113 100
rect 3121 94 3129 100
rect 3209 101 3237 114
rect 3209 94 3227 101
rect 2981 90 2985 94
rect 3089 90 3093 94
rect 3197 90 3201 94
rect 3305 90 3309 94
rect 3324 90 3328 94
rect 2969 86 2972 90
rect 2976 86 2980 90
rect 2984 86 2989 90
rect 2993 86 2998 90
rect 3002 86 3008 90
rect 3012 86 3016 90
rect 3020 86 3025 90
rect 3029 86 3034 90
rect 3038 86 3061 90
rect 3065 86 3070 90
rect 3074 86 3080 90
rect 3084 86 3088 90
rect 3092 86 3097 90
rect 3101 86 3106 90
rect 3110 86 3116 90
rect 3120 86 3124 90
rect 3128 86 3133 90
rect 3137 86 3142 90
rect 3146 86 3169 90
rect 3173 86 3178 90
rect 3182 86 3188 90
rect 3192 86 3196 90
rect 3200 86 3205 90
rect 3209 86 3214 90
rect 3218 86 3241 90
rect 3245 86 3250 90
rect 3254 86 3260 90
rect 3264 86 3268 90
rect 3272 86 3277 90
rect 3281 86 3286 90
rect 3290 86 3296 90
rect 3300 86 3304 90
rect 3308 86 3313 90
rect 3317 86 3323 90
rect 3327 86 3332 90
rect 3336 86 3341 90
rect 3345 87 3348 90
rect 3369 87 3373 318
rect 3345 86 3373 87
rect 2969 83 3373 86
rect 3058 74 3125 80
rect 3200 71 3206 72
rect 3272 71 3278 74
rect 3121 65 3278 71
rect 3305 63 3315 72
rect 2517 -215 2538 -211
rect 2545 -215 2554 -211
rect 2448 -221 2459 -216
rect 2525 -227 2529 -215
rect 2441 -237 2458 -227
rect 2470 -237 2529 -227
rect 2545 -220 2548 -215
rect 2561 -216 2759 -211
rect 2802 -118 3063 -113
rect 2561 -220 2564 -216
rect 2441 -244 2448 -237
rect 2536 -244 2540 -228
rect 2552 -244 2556 -228
rect 2441 -250 2574 -244
rect 2802 -259 2807 -118
rect 2968 -120 3063 -118
rect 2968 -124 2975 -120
rect 3056 -121 3063 -120
rect 2968 -131 2979 -124
rect 2953 -136 3345 -134
rect 2953 -140 2970 -136
rect 2974 -140 2979 -136
rect 2983 -140 2996 -136
rect 3000 -140 3006 -136
rect 3010 -140 3015 -136
rect 3019 -140 3032 -136
rect 3036 -140 3042 -136
rect 3046 -140 3051 -136
rect 3055 -140 3068 -136
rect 3072 -140 3078 -136
rect 3082 -140 3087 -136
rect 3091 -140 3104 -136
rect 3108 -140 3114 -136
rect 3118 -140 3123 -136
rect 3127 -140 3140 -136
rect 3144 -140 3150 -136
rect 3154 -140 3159 -136
rect 3163 -140 3176 -136
rect 3180 -140 3186 -136
rect 3190 -140 3195 -136
rect 3199 -140 3212 -136
rect 3216 -140 3222 -136
rect 3226 -140 3231 -136
rect 3235 -140 3248 -136
rect 3252 -140 3258 -136
rect 3262 -140 3267 -136
rect 3271 -140 3284 -136
rect 3288 -140 3294 -136
rect 3298 -140 3303 -136
rect 3307 -140 3320 -136
rect 3324 -140 3337 -136
rect 3341 -140 3345 -136
rect 2953 -142 3345 -140
rect 3061 -144 3065 -142
rect 3168 -144 3172 -142
rect 3136 -154 3160 -145
rect 3276 -144 3280 -142
rect 3244 -154 3268 -145
rect 3304 -144 3308 -142
rect 3321 -144 3325 -142
rect 3053 -167 3057 -154
rect 3124 -167 3128 -154
rect 3232 -167 3236 -154
rect 3312 -157 3316 -154
rect 3329 -155 3333 -154
rect 3312 -162 3321 -157
rect 3329 -160 3340 -155
rect 3312 -167 3316 -162
rect 3329 -167 3333 -160
rect 2992 -187 3016 -167
rect 3028 -181 3057 -167
rect 3028 -187 3048 -181
rect 3100 -181 3128 -167
rect 3100 -187 3112 -181
rect 3120 -187 3128 -181
rect 3208 -180 3236 -167
rect 3208 -187 3226 -180
rect 2980 -191 2984 -187
rect 3088 -191 3092 -187
rect 3196 -191 3200 -187
rect 3304 -191 3308 -187
rect 3321 -191 3325 -187
rect 2968 -195 2971 -191
rect 2975 -195 2979 -191
rect 2983 -195 2988 -191
rect 2992 -195 2997 -191
rect 3001 -195 3007 -191
rect 3011 -195 3015 -191
rect 3019 -195 3024 -191
rect 3028 -195 3033 -191
rect 3037 -195 3060 -191
rect 3064 -195 3069 -191
rect 3073 -195 3079 -191
rect 3083 -195 3087 -191
rect 3091 -195 3096 -191
rect 3100 -195 3105 -191
rect 3109 -195 3115 -191
rect 3119 -195 3123 -191
rect 3127 -195 3132 -191
rect 3136 -195 3141 -191
rect 3145 -195 3168 -191
rect 3172 -195 3177 -191
rect 3181 -195 3187 -191
rect 3191 -195 3195 -191
rect 3199 -195 3204 -191
rect 3208 -195 3213 -191
rect 3217 -195 3240 -191
rect 3244 -195 3249 -191
rect 3253 -195 3259 -191
rect 3263 -195 3267 -191
rect 3271 -195 3276 -191
rect 3280 -195 3285 -191
rect 3289 -195 3295 -191
rect 3299 -195 3303 -191
rect 3307 -195 3320 -191
rect 3324 -195 3329 -191
rect 3333 -195 3338 -191
rect 3342 -194 3345 -191
rect 3359 -194 3363 83
rect 3342 -195 3363 -194
rect 2968 -198 3363 -195
rect 3057 -207 3124 -201
rect 3199 -210 3205 -209
rect 3271 -210 3277 -207
rect 3120 -216 3277 -210
rect 3304 -218 3314 -209
rect 2562 -264 2807 -259
rect 2433 -389 2570 -386
rect 2433 -391 2532 -389
rect 2529 -393 2532 -391
rect 2536 -393 2545 -389
rect 2549 -393 2561 -389
rect 2565 -393 2570 -389
rect 2529 -394 2570 -393
rect 2536 -398 2540 -394
rect 2552 -398 2556 -394
rect 2448 -405 2467 -402
rect 2448 -406 2454 -405
rect 2465 -406 2467 -405
rect 2448 -426 2453 -406
rect 2457 -417 2462 -413
rect 2517 -414 2529 -410
rect 2462 -422 2467 -418
rect 2525 -426 2529 -414
rect 3121 -412 3278 -406
rect 3200 -413 3206 -412
rect 2544 -423 2548 -418
rect 2560 -423 2564 -418
rect 3058 -421 3125 -415
rect 3272 -415 3278 -412
rect 3305 -413 3315 -404
rect 2545 -426 2548 -423
rect 2561 -426 2564 -423
rect 3359 -424 3363 -198
rect 2517 -430 2538 -426
rect 2545 -430 2554 -426
rect 2448 -436 2459 -431
rect 2525 -442 2529 -430
rect 2441 -452 2458 -442
rect 2470 -452 2529 -442
rect 2545 -435 2548 -430
rect 2561 -431 2933 -426
rect 2969 -427 3363 -424
rect 2969 -431 2972 -427
rect 2976 -431 2980 -427
rect 2984 -431 2989 -427
rect 2993 -431 2998 -427
rect 3002 -431 3008 -427
rect 3012 -431 3016 -427
rect 3020 -431 3025 -427
rect 3029 -431 3034 -427
rect 3038 -431 3061 -427
rect 3065 -431 3070 -427
rect 3074 -431 3080 -427
rect 3084 -431 3088 -427
rect 3092 -431 3097 -427
rect 3101 -431 3106 -427
rect 3110 -431 3116 -427
rect 3120 -431 3124 -427
rect 3128 -431 3133 -427
rect 3137 -431 3142 -427
rect 3146 -431 3169 -427
rect 3173 -431 3178 -427
rect 3182 -431 3188 -427
rect 3192 -431 3196 -427
rect 3200 -431 3205 -427
rect 3209 -431 3214 -427
rect 3218 -431 3241 -427
rect 3245 -431 3250 -427
rect 3254 -431 3260 -427
rect 3264 -431 3268 -427
rect 3272 -431 3277 -427
rect 3281 -431 3286 -427
rect 3290 -431 3296 -427
rect 3300 -431 3304 -427
rect 3308 -431 3320 -427
rect 3324 -431 3329 -427
rect 3333 -428 3363 -427
rect 3333 -431 3343 -428
rect 2561 -435 2564 -431
rect 2441 -459 2448 -452
rect 2536 -459 2540 -443
rect 2552 -459 2556 -443
rect 2441 -462 2574 -459
rect 2412 -465 2574 -462
rect 2928 -494 2933 -431
rect 2981 -435 2985 -431
rect 3089 -435 3093 -431
rect 3197 -435 3201 -431
rect 3305 -435 3309 -431
rect 3321 -435 3325 -431
rect 2993 -455 3017 -435
rect 3029 -441 3049 -435
rect 3029 -455 3058 -441
rect 3101 -441 3113 -435
rect 3121 -441 3129 -435
rect 3101 -455 3129 -441
rect 3209 -442 3227 -435
rect 3209 -455 3237 -442
rect 3054 -468 3058 -455
rect 3125 -468 3129 -455
rect 3233 -468 3237 -455
rect 3313 -460 3317 -455
rect 3313 -465 3321 -460
rect 3329 -462 3333 -455
rect 3313 -468 3317 -465
rect 3329 -467 3340 -462
rect 3329 -468 3333 -467
rect 3137 -477 3161 -468
rect 3062 -480 3066 -478
rect 3245 -477 3269 -468
rect 3169 -480 3173 -478
rect 3277 -480 3281 -478
rect 3305 -480 3309 -478
rect 3321 -480 3325 -478
rect 2969 -482 3343 -480
rect 2969 -486 2971 -482
rect 2975 -486 2980 -482
rect 2984 -486 2997 -482
rect 3001 -486 3007 -482
rect 3011 -486 3016 -482
rect 3020 -486 3033 -482
rect 3037 -486 3043 -482
rect 3047 -486 3052 -482
rect 3056 -486 3069 -482
rect 3073 -486 3079 -482
rect 3083 -486 3088 -482
rect 3092 -486 3105 -482
rect 3109 -486 3115 -482
rect 3119 -486 3124 -482
rect 3128 -486 3141 -482
rect 3145 -486 3151 -482
rect 3155 -486 3160 -482
rect 3164 -486 3177 -482
rect 3181 -486 3187 -482
rect 3191 -486 3196 -482
rect 3200 -486 3213 -482
rect 3217 -486 3223 -482
rect 3227 -486 3232 -482
rect 3236 -486 3249 -482
rect 3253 -486 3259 -482
rect 3263 -486 3268 -482
rect 3272 -486 3285 -482
rect 3289 -486 3295 -482
rect 3299 -486 3304 -482
rect 3308 -486 3320 -482
rect 3324 -486 3337 -482
rect 3341 -486 3343 -482
rect 2969 -488 3343 -486
rect 2969 -494 2980 -491
rect 2928 -498 2980 -494
rect 2928 -499 2976 -498
rect 2969 -502 2976 -499
rect 3057 -502 3064 -501
rect 2969 -509 3064 -502
rect 3140 -543 3143 -488
rect 2013 -583 3064 -578
rect 1893 -590 1901 -585
rect 1893 -594 1895 -590
rect 1899 -594 1901 -590
rect 1893 -599 1901 -594
rect 1893 -603 1895 -599
rect 1899 -603 1901 -599
rect 1893 -609 1901 -603
rect 1893 -613 1895 -609
rect 1899 -613 1901 -609
rect 1893 -626 1901 -613
rect 1904 -617 1913 -593
rect 1950 -590 1957 -585
rect 1966 -590 1975 -584
rect 1954 -594 1957 -590
rect 1950 -598 1957 -594
rect 1954 -602 1957 -598
rect 1950 -608 1957 -602
rect 1954 -612 1957 -608
rect 1950 -617 1957 -612
rect 1954 -621 1957 -617
rect 1741 -635 1754 -629
rect 1734 -653 1754 -635
rect 1779 -630 1781 -626
rect 1785 -630 1787 -626
rect 1779 -635 1787 -630
rect 1779 -639 1781 -635
rect 1785 -639 1787 -635
rect 1779 -645 1787 -639
rect 1779 -649 1781 -645
rect 1785 -649 1787 -645
rect 1723 -661 1730 -657
rect 1723 -662 1734 -661
rect 1705 -741 1711 -662
rect 1723 -666 1726 -662
rect 1730 -665 1734 -662
rect 1779 -662 1787 -649
rect 1723 -670 1730 -666
rect 1723 -674 1726 -670
rect 1723 -680 1730 -674
rect 1723 -684 1726 -680
rect 1723 -689 1730 -684
rect 1779 -666 1781 -662
rect 1785 -666 1787 -662
rect 1779 -671 1787 -666
rect 1779 -675 1781 -671
rect 1785 -675 1787 -671
rect 1779 -681 1787 -675
rect 1779 -685 1781 -681
rect 1785 -685 1787 -681
rect 1779 -689 1787 -685
rect 1723 -693 1726 -689
rect 1777 -693 1787 -689
rect 1893 -630 1895 -626
rect 1899 -630 1901 -626
rect 1913 -629 1939 -625
rect 1893 -635 1901 -630
rect 1893 -639 1895 -635
rect 1899 -639 1901 -635
rect 1893 -645 1901 -639
rect 1893 -649 1895 -645
rect 1899 -649 1901 -645
rect 1893 -662 1901 -649
rect 1926 -635 1939 -629
rect 1926 -653 1946 -635
rect 1950 -644 1957 -621
rect 1954 -648 1957 -644
rect 1950 -653 1957 -648
rect 1954 -657 1957 -653
rect 1969 -656 1975 -590
rect 2969 -585 3064 -583
rect 2969 -589 2976 -585
rect 3057 -586 3064 -585
rect 2969 -596 2980 -589
rect 3140 -599 3143 -548
rect 2969 -601 3342 -599
rect 2969 -605 2971 -601
rect 2975 -605 2980 -601
rect 2984 -605 2997 -601
rect 3001 -605 3007 -601
rect 3011 -605 3016 -601
rect 3020 -605 3033 -601
rect 3037 -605 3043 -601
rect 3047 -605 3052 -601
rect 3056 -605 3069 -601
rect 3073 -605 3079 -601
rect 3083 -605 3088 -601
rect 3092 -605 3105 -601
rect 3109 -605 3115 -601
rect 3119 -605 3124 -601
rect 3128 -605 3141 -601
rect 3145 -605 3151 -601
rect 3155 -605 3160 -601
rect 3164 -605 3177 -601
rect 3181 -605 3187 -601
rect 3191 -605 3196 -601
rect 3200 -605 3213 -601
rect 3217 -605 3223 -601
rect 3227 -605 3232 -601
rect 3236 -605 3249 -601
rect 3253 -605 3259 -601
rect 3263 -605 3268 -601
rect 3272 -605 3285 -601
rect 3289 -605 3295 -601
rect 3299 -605 3304 -601
rect 3308 -605 3320 -601
rect 3324 -605 3337 -601
rect 3341 -605 3342 -601
rect 2969 -607 3342 -605
rect 3062 -609 3066 -607
rect 3169 -609 3173 -607
rect 3137 -619 3161 -610
rect 3277 -609 3281 -607
rect 3245 -619 3269 -610
rect 3305 -609 3309 -607
rect 3321 -609 3325 -607
rect 3054 -632 3058 -619
rect 3125 -632 3129 -619
rect 3233 -632 3237 -619
rect 3313 -622 3317 -619
rect 3329 -620 3333 -619
rect 3313 -627 3321 -622
rect 3329 -625 3341 -620
rect 3313 -632 3317 -627
rect 3329 -632 3333 -625
rect 2993 -652 3017 -632
rect 3029 -646 3058 -632
rect 3029 -652 3049 -646
rect 3101 -646 3129 -632
rect 3101 -652 3113 -646
rect 3121 -652 3129 -646
rect 3209 -645 3237 -632
rect 3209 -652 3227 -645
rect 2981 -656 2985 -652
rect 3089 -656 3093 -652
rect 3197 -656 3201 -652
rect 3305 -656 3309 -652
rect 3321 -656 3325 -652
rect 1950 -661 1957 -657
rect 1893 -666 1895 -662
rect 1899 -666 1901 -662
rect 1946 -662 1957 -661
rect 1968 -662 1975 -656
rect 1946 -665 1950 -662
rect 1893 -671 1901 -666
rect 1893 -675 1895 -671
rect 1899 -675 1901 -671
rect 1893 -681 1901 -675
rect 1893 -685 1895 -681
rect 1899 -685 1901 -681
rect 1893 -689 1901 -685
rect 1954 -666 1957 -662
rect 1950 -670 1957 -666
rect 1954 -674 1957 -670
rect 1950 -680 1957 -674
rect 1954 -684 1957 -680
rect 1950 -689 1957 -684
rect 1723 -716 1730 -693
rect 1723 -720 1726 -716
rect 1723 -725 1730 -720
rect 1723 -729 1726 -725
rect 1767 -725 1776 -701
rect 1779 -698 1787 -693
rect 1893 -693 1903 -689
rect 1954 -693 1957 -689
rect 1893 -698 1901 -693
rect 1779 -702 1781 -698
rect 1785 -702 1787 -698
rect 1779 -707 1787 -702
rect 1779 -711 1781 -707
rect 1785 -711 1787 -707
rect 1779 -715 1787 -711
rect 1893 -702 1895 -698
rect 1899 -702 1901 -698
rect 1893 -707 1901 -702
rect 1893 -711 1895 -707
rect 1899 -711 1901 -707
rect 1893 -715 1901 -711
rect 1779 -717 1838 -715
rect 1779 -721 1781 -717
rect 1785 -720 1838 -717
rect 1843 -717 1901 -715
rect 1843 -720 1895 -717
rect 1785 -721 1787 -720
rect 1714 -804 1720 -737
rect 1723 -734 1730 -729
rect 1723 -738 1726 -734
rect 1723 -742 1730 -738
rect 1723 -746 1726 -742
rect 1723 -752 1730 -746
rect 1723 -756 1726 -752
rect 1723 -761 1730 -756
rect 1723 -765 1726 -761
rect 1734 -737 1767 -733
rect 1779 -734 1787 -721
rect 1734 -741 1754 -737
rect 1740 -749 1754 -741
rect 1734 -761 1754 -749
rect 1779 -738 1781 -734
rect 1785 -738 1787 -734
rect 1779 -743 1787 -738
rect 1779 -747 1781 -743
rect 1785 -747 1787 -743
rect 1779 -753 1787 -747
rect 1779 -757 1781 -753
rect 1785 -757 1787 -753
rect 1723 -769 1730 -765
rect 1723 -770 1734 -769
rect 1723 -774 1726 -770
rect 1730 -773 1734 -770
rect 1779 -770 1787 -757
rect 1893 -721 1895 -720
rect 1899 -721 1901 -717
rect 1893 -734 1901 -721
rect 1904 -725 1913 -701
rect 1950 -716 1957 -693
rect 1954 -720 1957 -716
rect 1950 -725 1957 -720
rect 1954 -729 1957 -725
rect 1893 -738 1895 -734
rect 1899 -738 1901 -734
rect 1913 -737 1946 -733
rect 1893 -743 1901 -738
rect 1893 -747 1895 -743
rect 1899 -747 1901 -743
rect 1893 -753 1901 -747
rect 1893 -757 1895 -753
rect 1899 -757 1901 -753
rect 1893 -770 1901 -757
rect 1926 -741 1946 -737
rect 1926 -749 1940 -741
rect 1926 -761 1946 -749
rect 1950 -734 1957 -729
rect 1954 -738 1957 -734
rect 1950 -742 1957 -738
rect 1954 -746 1957 -742
rect 1950 -752 1957 -746
rect 1954 -756 1957 -752
rect 1950 -761 1957 -756
rect 1954 -765 1957 -761
rect 1950 -769 1957 -765
rect 1723 -778 1730 -774
rect 1723 -782 1726 -778
rect 1723 -788 1730 -782
rect 1723 -792 1726 -788
rect 1723 -797 1730 -792
rect 1779 -774 1781 -770
rect 1785 -774 1787 -770
rect 1779 -779 1787 -774
rect 1779 -783 1781 -779
rect 1785 -783 1787 -779
rect 1779 -789 1787 -783
rect 1779 -793 1781 -789
rect 1785 -793 1787 -789
rect 1779 -796 1787 -793
rect 1723 -801 1726 -797
rect 1777 -800 1787 -796
rect 1893 -774 1895 -770
rect 1899 -774 1901 -770
rect 1946 -770 1957 -769
rect 1946 -773 1950 -770
rect 1893 -779 1901 -774
rect 1893 -783 1895 -779
rect 1899 -783 1901 -779
rect 1893 -789 1901 -783
rect 1893 -793 1895 -789
rect 1899 -793 1901 -789
rect 1893 -796 1901 -793
rect 1954 -774 1957 -770
rect 1950 -778 1957 -774
rect 1954 -782 1957 -778
rect 1950 -788 1957 -782
rect 1954 -792 1957 -788
rect 1723 -824 1730 -801
rect 1723 -828 1726 -824
rect 1723 -833 1730 -828
rect 1723 -837 1726 -833
rect 1740 -808 1767 -804
rect 1779 -806 1787 -800
rect 1800 -805 1808 -798
rect 1740 -813 1754 -808
rect 1734 -833 1754 -813
rect 1779 -810 1781 -806
rect 1785 -810 1787 -806
rect 1779 -815 1787 -810
rect 1779 -819 1781 -815
rect 1785 -819 1787 -815
rect 1779 -825 1787 -819
rect 1779 -829 1781 -825
rect 1785 -829 1787 -825
rect 1723 -842 1730 -837
rect 1723 -846 1726 -842
rect 1723 -850 1730 -846
rect 1723 -854 1726 -850
rect 1723 -860 1730 -854
rect 1723 -864 1726 -860
rect 1723 -869 1730 -864
rect 1723 -873 1726 -869
rect 1734 -869 1754 -845
rect 1779 -842 1787 -829
rect 1779 -846 1781 -842
rect 1785 -846 1787 -842
rect 1779 -851 1787 -846
rect 1779 -855 1781 -851
rect 1785 -855 1787 -851
rect 1779 -861 1787 -855
rect 1779 -865 1781 -861
rect 1785 -865 1787 -861
rect 1723 -877 1730 -873
rect 1723 -878 1734 -877
rect 1723 -882 1726 -878
rect 1730 -881 1734 -878
rect 1779 -878 1787 -865
rect 1723 -886 1730 -882
rect 1723 -890 1726 -886
rect 1723 -893 1730 -890
rect 1779 -882 1781 -878
rect 1785 -882 1787 -878
rect 1779 -887 1787 -882
rect 1779 -891 1781 -887
rect 1785 -891 1787 -887
rect 1779 -893 1787 -891
rect 1790 -886 1797 -882
rect 1801 -886 1808 -805
rect 1790 -893 1808 -886
rect 1872 -805 1880 -798
rect 1893 -800 1903 -796
rect 1950 -797 1957 -792
rect 1872 -886 1879 -805
rect 1893 -806 1901 -800
rect 1954 -801 1957 -797
rect 1893 -810 1895 -806
rect 1899 -810 1901 -806
rect 1913 -808 1940 -804
rect 1893 -815 1901 -810
rect 1893 -819 1895 -815
rect 1899 -819 1901 -815
rect 1893 -825 1901 -819
rect 1893 -829 1895 -825
rect 1899 -829 1901 -825
rect 1893 -842 1901 -829
rect 1926 -813 1940 -808
rect 1926 -833 1946 -813
rect 1950 -824 1957 -801
rect 1960 -804 1966 -737
rect 1969 -741 1975 -662
rect 2969 -660 2972 -656
rect 2976 -660 2980 -656
rect 2984 -660 2989 -656
rect 2993 -660 2998 -656
rect 3002 -660 3008 -656
rect 3012 -660 3016 -656
rect 3020 -660 3025 -656
rect 3029 -660 3034 -656
rect 3038 -660 3061 -656
rect 3065 -660 3070 -656
rect 3074 -660 3080 -656
rect 3084 -660 3088 -656
rect 3092 -660 3097 -656
rect 3101 -660 3106 -656
rect 3110 -660 3116 -656
rect 3120 -660 3124 -656
rect 3128 -660 3133 -656
rect 3137 -660 3142 -656
rect 3146 -660 3169 -656
rect 3173 -660 3178 -656
rect 3182 -660 3188 -656
rect 3192 -660 3196 -656
rect 3200 -660 3205 -656
rect 3209 -660 3214 -656
rect 3218 -660 3241 -656
rect 3245 -660 3250 -656
rect 3254 -660 3260 -656
rect 3264 -660 3268 -656
rect 3272 -660 3277 -656
rect 3281 -660 3286 -656
rect 3290 -660 3296 -656
rect 3300 -660 3304 -656
rect 3308 -660 3320 -656
rect 3324 -660 3329 -656
rect 3333 -659 3342 -656
rect 3359 -659 3363 -428
rect 3333 -660 3363 -659
rect 2969 -663 3363 -660
rect 3058 -672 3125 -666
rect 3200 -675 3206 -674
rect 3272 -675 3278 -672
rect 3121 -681 3278 -675
rect 3305 -683 3315 -674
rect 1954 -828 1957 -824
rect 1950 -833 1957 -828
rect 1954 -837 1957 -833
rect 1893 -846 1895 -842
rect 1899 -846 1901 -842
rect 1893 -851 1901 -846
rect 1893 -855 1895 -851
rect 1899 -855 1901 -851
rect 1893 -861 1901 -855
rect 1893 -865 1895 -861
rect 1899 -865 1901 -861
rect 1883 -886 1890 -882
rect 1872 -893 1890 -886
rect 1893 -878 1901 -865
rect 1926 -869 1946 -845
rect 1950 -842 1957 -837
rect 1954 -846 1957 -842
rect 1950 -850 1957 -846
rect 1954 -854 1957 -850
rect 1950 -860 1957 -854
rect 1954 -864 1957 -860
rect 1950 -869 1957 -864
rect 1954 -873 1957 -869
rect 1950 -877 1957 -873
rect 1893 -882 1895 -878
rect 1899 -882 1901 -878
rect 1946 -878 1957 -877
rect 1946 -881 1950 -878
rect 1893 -887 1901 -882
rect 1893 -891 1895 -887
rect 1899 -891 1901 -887
rect 1893 -893 1901 -891
rect 1954 -882 1957 -878
rect 1950 -886 1957 -882
rect 1954 -890 1957 -886
rect 1950 -893 1957 -890
rect 1723 -905 1727 -893
rect 1953 -905 1957 -893
rect 3359 -905 3363 -663
rect 1169 -909 3363 -905
<< m2contact >>
rect 1736 430 1742 439
rect 1727 367 1733 375
rect 1756 430 1762 439
rect 1962 430 1968 439
rect 1756 367 1762 375
rect 1858 375 1863 380
rect 1962 367 1968 375
rect 1982 430 1988 439
rect 1991 367 1997 375
rect 1756 251 1763 261
rect 3305 342 3315 349
rect 3113 334 3121 340
rect 3049 325 3058 331
rect 3049 305 3058 311
rect 3113 305 3121 311
rect 3227 304 3237 311
rect 1718 173 1725 183
rect 1529 147 1539 154
rect 1337 139 1345 145
rect 1273 130 1282 136
rect 1273 110 1282 116
rect 1337 110 1345 116
rect 1451 109 1461 116
rect 1330 15 1335 20
rect 1961 251 1968 261
rect 1999 173 2006 183
rect 1939 40 1944 45
rect 1781 31 1786 36
rect 1761 4 1766 9
rect 1659 -55 1664 -50
rect 1273 -83 1282 -77
rect 1337 -83 1345 -77
rect 1451 -83 1461 -76
rect 1273 -103 1282 -97
rect 1337 -112 1345 -106
rect 1529 -121 1539 -114
rect 1731 -30 1736 -25
rect 1722 -39 1727 -34
rect 1524 -274 1534 -267
rect 1332 -282 1340 -276
rect 1268 -291 1277 -285
rect 1268 -311 1277 -305
rect 1332 -311 1340 -305
rect 1446 -312 1456 -305
rect 1677 -336 1682 -331
rect 1698 -156 1704 -151
rect 1819 -30 1824 -25
rect 1810 -39 1815 -34
rect 1764 -156 1770 -151
rect 1908 -30 1913 -25
rect 1899 -39 1904 -34
rect 1852 -156 1858 -151
rect 1941 -156 1947 -151
rect 1996 -30 2001 -25
rect 1987 -39 1992 -34
rect 2073 -96 2078 -91
rect 1966 -156 1971 -151
rect 2242 -65 2247 -60
rect 2262 -103 2267 -98
rect 2029 -156 2035 -151
rect 2403 -30 2408 -25
rect 2344 -157 2349 -152
rect 2381 -168 2386 -163
rect 2006 -194 2011 -189
rect 2085 -194 2090 -189
rect 2235 -194 2240 -189
rect 2365 -194 2370 -189
rect 2015 -202 2020 -197
rect 2457 -21 2462 -16
rect 3183 204 3188 209
rect 2448 -30 2453 -25
rect 2574 -64 2579 -58
rect 2025 -210 2030 -205
rect 2184 -210 2189 -205
rect 2334 -210 2339 -205
rect 2403 -210 2408 -205
rect 2085 -231 2090 -226
rect 2290 -247 2295 -242
rect 2172 -255 2177 -250
rect 2064 -263 2069 -258
rect 2161 -271 2166 -266
rect 2325 -271 2330 -266
rect 2075 -287 2080 -282
rect 2244 -287 2249 -282
rect 1959 -295 1964 -290
rect 1913 -329 1918 -324
rect 1394 -413 1399 -408
rect 1674 -380 1679 -375
rect 1811 -397 1816 -392
rect 1758 -416 1763 -411
rect 1268 -517 1277 -511
rect 1332 -517 1340 -511
rect 1446 -517 1456 -510
rect 1268 -537 1277 -531
rect 1332 -546 1340 -540
rect 1524 -555 1534 -548
rect 1696 -557 1703 -547
rect 1734 -635 1741 -625
rect 2262 -396 2267 -391
rect 2343 -407 2348 -402
rect 1977 -557 1984 -547
rect 2457 -207 2462 -202
rect 3049 94 3058 100
rect 3113 94 3121 100
rect 3227 94 3237 101
rect 3049 74 3058 80
rect 3113 65 3121 71
rect 3305 56 3315 63
rect 2448 -216 2453 -211
rect 2574 -250 2579 -244
rect 2945 -142 2953 -134
rect 3048 -187 3057 -181
rect 3112 -187 3120 -181
rect 3226 -187 3236 -180
rect 3048 -207 3057 -201
rect 3112 -216 3120 -210
rect 3304 -225 3314 -218
rect 2557 -264 2562 -259
rect 2457 -422 2462 -417
rect 3305 -404 3315 -397
rect 3113 -412 3121 -406
rect 3049 -421 3058 -415
rect 2448 -431 2453 -426
rect 2574 -465 2579 -459
rect 3049 -441 3058 -435
rect 3113 -441 3121 -435
rect 3227 -442 3237 -435
rect 3138 -548 3143 -543
rect 1939 -635 1946 -625
rect 3049 -652 3058 -646
rect 3113 -652 3121 -646
rect 3227 -652 3237 -645
rect 1838 -720 1843 -715
rect 1705 -749 1711 -741
rect 1714 -813 1720 -804
rect 1734 -749 1740 -741
rect 1940 -749 1946 -741
rect 1734 -813 1740 -804
rect 1940 -813 1946 -804
rect 3049 -672 3058 -666
rect 3113 -681 3121 -675
rect 3305 -690 3315 -683
rect 1969 -749 1975 -741
rect 1960 -813 1966 -804
<< pm12contact >>
rect 1812 465 1819 472
rect 1905 465 1912 472
rect 1815 390 1821 396
rect 1903 390 1909 396
rect 1813 318 1819 324
rect 1905 318 1911 324
rect 1813 246 1819 252
rect 1905 246 1911 252
rect 1240 53 1247 60
rect 1316 51 1322 57
rect 1388 53 1394 59
rect 1460 53 1466 59
rect 1240 -27 1247 -20
rect 1316 -24 1322 -18
rect 3016 248 3023 255
rect 3092 246 3098 252
rect 3164 248 3170 254
rect 1388 -26 1394 -20
rect 1460 -26 1466 -20
rect 1235 -368 1242 -361
rect 1311 -370 1317 -364
rect 1383 -368 1389 -362
rect 2064 -104 2069 -99
rect 2075 -133 2080 -128
rect 2085 -145 2090 -140
rect 2172 -43 2177 -38
rect 2184 -55 2189 -50
rect 2284 -82 2289 -77
rect 2161 -133 2166 -128
rect 2244 -121 2249 -116
rect 2235 -133 2240 -128
rect 2334 -121 2339 -116
rect 2325 -133 2330 -128
rect 3236 248 3242 254
rect 2025 -314 2030 -309
rect 2015 -339 2020 -334
rect 2006 -350 2011 -345
rect 1455 -368 1461 -362
rect 1699 -371 1704 -366
rect 1714 -372 1719 -367
rect 1758 -371 1763 -366
rect 1770 -371 1775 -366
rect 1811 -371 1816 -366
rect 1822 -371 1827 -366
rect 1866 -371 1871 -366
rect 1878 -371 1883 -366
rect 1235 -461 1242 -454
rect 1311 -458 1317 -452
rect 1383 -460 1389 -454
rect 1455 -460 1461 -454
rect 2078 -370 2083 -365
rect 3016 150 3023 157
rect 3092 153 3098 159
rect 3164 151 3170 157
rect 3236 151 3242 157
rect 3015 -131 3022 -124
rect 3091 -128 3097 -122
rect 3163 -130 3169 -124
rect 3235 -130 3241 -124
rect 3016 -498 3023 -491
rect 3092 -500 3098 -494
rect 3164 -498 3170 -492
rect 3236 -498 3242 -492
rect 1791 -626 1797 -620
rect 1883 -626 1889 -620
rect 3016 -596 3023 -589
rect 3092 -593 3098 -587
rect 3164 -595 3170 -589
rect 3236 -595 3242 -589
rect 1791 -698 1797 -692
rect 1883 -698 1889 -692
rect 1793 -770 1799 -764
rect 1881 -770 1887 -764
rect 1790 -846 1797 -839
rect 1883 -846 1890 -839
<< ndm12contact >>
rect 1697 -295 1702 -290
rect 1733 -315 1738 -310
rect 1753 -295 1758 -290
rect 1789 -316 1794 -311
rect 1806 -295 1811 -290
rect 1841 -316 1846 -311
rect 1862 -295 1867 -290
rect 1897 -316 1902 -311
rect 1917 -316 1922 -311
rect 1935 -316 1940 -311
<< metal2 >>
rect 1129 595 3532 599
rect 1129 27 1134 595
rect 1857 593 3532 595
rect 1857 479 1862 593
rect 1812 474 1912 479
rect 1812 472 1841 474
rect 1742 430 1756 439
rect 1835 396 1841 472
rect 1821 390 1841 396
rect 1733 367 1756 375
rect 1835 324 1841 390
rect 1883 472 1912 474
rect 1883 396 1889 472
rect 1968 430 1982 439
rect 1883 390 1903 396
rect 1819 318 1841 324
rect 1718 251 1756 261
rect 1835 252 1841 318
rect 1718 183 1725 251
rect 1819 246 1841 252
rect 1451 147 1529 154
rect 1273 116 1282 130
rect 1337 116 1345 139
rect 1451 116 1461 147
rect 1858 110 1863 375
rect 1883 324 1889 390
rect 1968 367 1991 375
rect 3227 342 3305 349
rect 1883 318 1905 324
rect 1883 252 1889 318
rect 3049 311 3058 325
rect 3113 311 3121 334
rect 3227 311 3237 342
rect 1883 246 1905 252
rect 1968 251 2006 261
rect 1999 183 2006 251
rect 3009 232 3016 255
rect 3092 232 3098 246
rect 3164 232 3170 248
rect 3236 232 3242 248
rect 3009 226 3242 232
rect 2880 204 3183 209
rect 2880 110 2885 204
rect 3235 199 3242 226
rect 3526 199 3532 593
rect 3235 194 3532 199
rect 3235 178 3242 194
rect 3009 173 3242 178
rect 3009 150 3016 173
rect 3092 159 3098 173
rect 3164 157 3170 173
rect 3236 157 3242 173
rect 1595 105 2885 110
rect 1233 37 1240 60
rect 1316 37 1322 51
rect 1388 37 1394 53
rect 1460 37 1466 53
rect 1233 31 1466 37
rect 1233 27 1238 31
rect 1129 22 1238 27
rect 1129 -401 1134 22
rect 1233 2 1238 22
rect 1595 20 1600 105
rect 1335 15 1600 20
rect 1233 -4 1466 2
rect 1233 -27 1240 -4
rect 1316 -18 1322 -4
rect 1388 -20 1394 -4
rect 1460 -20 1466 -4
rect 1273 -97 1282 -83
rect 1337 -106 1345 -83
rect 1451 -114 1461 -83
rect 1451 -121 1529 -114
rect 1446 -274 1524 -267
rect 1268 -305 1277 -291
rect 1332 -305 1340 -282
rect 1446 -305 1456 -274
rect 1228 -384 1235 -361
rect 1311 -384 1317 -370
rect 1383 -384 1389 -368
rect 1455 -384 1461 -368
rect 1228 -390 1461 -384
rect 1228 -401 1233 -390
rect 1129 -407 1233 -401
rect 1129 -921 1134 -407
rect 1228 -432 1233 -407
rect 1595 -408 1600 15
rect 1399 -413 1600 -408
rect 1228 -438 1461 -432
rect 1228 -461 1235 -438
rect 1311 -452 1317 -438
rect 1383 -454 1389 -438
rect 1455 -454 1461 -438
rect 1595 -453 1600 -413
rect 1614 40 1939 45
rect 1944 40 2001 45
rect 1614 -429 1619 40
rect 1623 31 1781 36
rect 1786 31 1992 36
rect 1623 -420 1628 31
rect 1632 22 1913 27
rect 1632 -411 1637 22
rect 1641 13 1904 18
rect 1641 -402 1646 13
rect 1650 4 1761 9
rect 1766 4 1824 9
rect 1650 -393 1655 4
rect 1659 -5 1815 0
rect 1659 -50 1664 -5
rect 1659 -384 1664 -55
rect 1668 -14 1736 -9
rect 1668 -375 1673 -14
rect 1677 -24 1727 -18
rect 1677 -331 1682 -24
rect 1722 -34 1727 -24
rect 1731 -25 1736 -14
rect 1810 -34 1815 -5
rect 1819 -25 1824 4
rect 1899 -34 1904 13
rect 1908 -25 1913 22
rect 1987 -34 1992 31
rect 1996 -25 2001 40
rect 2073 1 2409 6
rect 2073 -91 2078 1
rect 2404 -16 2409 1
rect 2404 -21 2457 -16
rect 2408 -30 2448 -25
rect 1704 -156 1764 -151
rect 1770 -156 1852 -151
rect 1858 -156 1941 -151
rect 1947 -156 1966 -151
rect 1971 -156 2029 -151
rect 1698 -290 1702 -156
rect 1966 -157 1971 -156
rect 1702 -295 1753 -290
rect 1758 -295 1806 -290
rect 1811 -295 1862 -290
rect 1867 -295 1959 -290
rect 1733 -310 1738 -295
rect 1789 -311 1794 -295
rect 1841 -311 1846 -295
rect 1897 -311 1902 -295
rect 1917 -311 1922 -295
rect 1935 -311 1940 -295
rect 1677 -366 1682 -336
rect 1677 -371 1699 -366
rect 1714 -375 1719 -372
rect 1668 -380 1674 -375
rect 1679 -380 1719 -375
rect 1758 -384 1763 -371
rect 1659 -389 1763 -384
rect 1770 -393 1775 -371
rect 1650 -398 1775 -393
rect 1811 -392 1816 -371
rect 1811 -402 1816 -397
rect 1641 -407 1816 -402
rect 1822 -411 1827 -371
rect 1632 -416 1758 -411
rect 1763 -416 1827 -411
rect 1866 -420 1871 -371
rect 1623 -425 1871 -420
rect 1878 -429 1883 -371
rect 1614 -434 1883 -429
rect 1913 -426 1918 -329
rect 2006 -345 2011 -194
rect 2015 -334 2020 -202
rect 2025 -309 2030 -210
rect 2064 -258 2069 -104
rect 2075 -282 2080 -133
rect 2085 -189 2090 -145
rect 2085 -365 2090 -231
rect 2161 -266 2166 -133
rect 2172 -250 2177 -43
rect 2184 -205 2189 -55
rect 2242 -68 2247 -65
rect 2242 -73 2433 -68
rect 2289 -82 2295 -77
rect 2235 -189 2240 -133
rect 2244 -282 2249 -121
rect 2083 -370 2090 -365
rect 2262 -391 2267 -103
rect 2290 -242 2295 -82
rect 2325 -266 2330 -133
rect 2334 -205 2339 -121
rect 2344 -402 2348 -157
rect 2365 -417 2370 -194
rect 2381 -259 2386 -168
rect 2428 -202 2433 -73
rect 2428 -207 2457 -202
rect 2403 -211 2408 -210
rect 2403 -216 2448 -211
rect 2574 -244 2579 -64
rect 2381 -264 2557 -259
rect 2574 -314 2579 -250
rect 2880 -135 2885 105
rect 3049 80 3058 94
rect 3113 71 3121 94
rect 3227 63 3237 94
rect 3227 56 3305 63
rect 3526 -107 3532 194
rect 3008 -111 3532 -107
rect 3008 -131 3015 -111
rect 3091 -122 3097 -111
rect 3163 -124 3169 -111
rect 3235 -124 3241 -111
rect 2880 -142 2945 -135
rect 2880 -314 2885 -142
rect 3048 -201 3057 -187
rect 3112 -210 3120 -187
rect 3226 -218 3236 -187
rect 3226 -225 3304 -218
rect 2574 -319 2885 -314
rect 2365 -422 2457 -417
rect 1913 -431 2448 -426
rect 1595 -458 1843 -453
rect 1268 -531 1277 -517
rect 1332 -540 1340 -517
rect 1446 -548 1456 -517
rect 1446 -555 1524 -548
rect 1696 -625 1703 -557
rect 1696 -635 1734 -625
rect 1797 -626 1819 -620
rect 1813 -692 1819 -626
rect 1797 -698 1819 -692
rect 1711 -749 1734 -741
rect 1813 -764 1819 -698
rect 1838 -715 1843 -458
rect 2574 -459 2579 -319
rect 2880 -543 2885 -319
rect 3227 -404 3305 -397
rect 3049 -435 3058 -421
rect 3113 -435 3121 -412
rect 3227 -435 3237 -404
rect 3009 -514 3016 -491
rect 3092 -514 3098 -500
rect 3164 -514 3170 -498
rect 3236 -514 3242 -498
rect 3009 -519 3242 -514
rect 2880 -548 3138 -543
rect 3235 -544 3242 -519
rect 3526 -544 3532 -111
rect 1861 -626 1883 -620
rect 1977 -625 1984 -557
rect 3235 -549 3532 -544
rect 3235 -567 3242 -549
rect 3009 -573 3242 -567
rect 3009 -596 3016 -573
rect 3092 -587 3098 -573
rect 3164 -589 3170 -573
rect 3236 -589 3242 -573
rect 1861 -692 1867 -626
rect 1946 -635 1984 -625
rect 3049 -666 3058 -652
rect 3113 -675 3121 -652
rect 3227 -683 3237 -652
rect 3227 -690 3305 -683
rect 1861 -698 1883 -692
rect 1799 -770 1819 -764
rect 1720 -813 1734 -804
rect 1813 -846 1819 -770
rect 1790 -848 1819 -846
rect 1861 -764 1867 -698
rect 1946 -749 1969 -741
rect 1861 -770 1881 -764
rect 1861 -846 1867 -770
rect 1946 -813 1960 -804
rect 1861 -848 1890 -846
rect 1790 -853 1890 -848
rect 1839 -920 1844 -853
rect 3526 -920 3532 -549
rect 1839 -921 3532 -920
rect 1129 -924 3532 -921
rect 1129 -925 3531 -924
rect 1129 -926 1844 -925
<< labels >>
rlabel metal1 1776 -12 1776 -12 1 vdd
rlabel metal1 1767 -115 1767 -115 1 gnd
rlabel m2contact 1915 -326 1915 -326 1 C1
rlabel metal1 2088 -119 2088 -119 1 1
rlabel metal1 2164 -124 2164 -124 1 2
rlabel metal1 2239 -110 2239 -110 1 3
rlabel metal1 2239 -62 2239 -62 1 C3
rlabel metal1 2334 -111 2334 -111 1 5
rlabel metal1 2251 -34 2251 -34 1 4
rlabel metal1 2017 -356 2017 -356 1 6
rlabel metal1 2014 -409 2014 -409 1 C4
rlabel metal1 2073 -95 2073 -95 1 C2
rlabel metal1 2562 -429 2562 -429 1 S02
rlabel metal1 2562 -28 2562 -28 1 S03
rlabel metal1 2562 -214 2562 -214 1 S04
rlabel metal1 1803 -876 1803 -876 1 b02
rlabel metal1 1874 -874 1874 -874 1 a02
rlabel metal1 1827 502 1827 502 1 a01
rlabel metal1 1896 499 1896 499 1 b01
rlabel metal1 1215 45 1215 45 1 b03
rlabel metal1 1208 -13 1208 -13 1 a03
rlabel metal1 1209 -376 1209 -376 1 a04
rlabel metal1 1209 -445 1209 -445 1 b04
rlabel metal1 3321 284 3321 284 1 S3
rlabel metal1 3318 122 3318 122 1 S4
rlabel metal1 3319 -160 3319 -160 1 S1
rlabel metal1 3320 -463 3320 -463 1 S2
rlabel polycontact 3323 -625 3323 -625 1 S5
rlabel metal2 3528 -187 3528 -187 7 clk
rlabel metal2 1999 -2 1999 -2 1 b1
rlabel metal2 1990 -1 1990 -1 1 a1
rlabel metal2 1911 -2 1911 -2 1 b2
rlabel metal2 1901 -1 1901 -1 1 a2
rlabel metal2 1822 -2 1822 -2 1 b3
rlabel metal2 1806 -2 1806 -2 1 a3
rlabel metal2 1703 -23 1703 -23 1 a4
rlabel metal2 1669 -23 1669 -23 1 b4
rlabel metal1 1998 -140 1998 -140 1 p0
rlabel metal1 1909 -140 1909 -140 1 p1
rlabel metal1 1822 -139 1822 -139 1 p2
rlabel metal1 1729 -140 1729 -140 1 p3
rlabel metal1 2031 -228 2031 -228 1 1g3
rlabel metal1 2033 -237 2033 -237 1 g3
rlabel metal1 2035 -245 2035 -245 1 1g2
rlabel metal1 2039 -253 2039 -253 1 g2
rlabel metal1 2041 -261 2041 -261 1 1g1
rlabel metal1 2041 -268 2041 -268 1 g1
rlabel metal1 1946 -325 1946 -325 1 g0
rlabel metal1 1892 -329 1892 -329 1 1g0
<< end >>
